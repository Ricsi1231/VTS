��   K�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_  �$$C�LASS  ������D��D�VERSION�  ���/IRTUA�L-9LOOR� G��DD<x$p?�������k,  1 <DwX< y�����D'����	/��Z�Zm//��/_/�/�/�/$ ��/�/	?';�$M�NU>A\"� 
 <��4/d?��[? }?�?�?�?�?�?�?O`�?O1O_OEI cO �OwO�O�O�O�O�O_��O_E_�;5NUM  �����92�TOOLC?\ �
Y;�]2��F%4�P�RQ�d���F4�PSQ?�唊Aa��C���GOY_	oAOo ?o%o7oYo�omo�o�o 1_�o�o�o�o;! CqWy���� ��Z�Vy�Wy