��   ��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����BIN_CFG�_TX 	$E�NTRIES  $Q0FP?UNG1F1O2F�2OPz ?CNE�TG���DHC�P_CTRL. � 0 7 AB�LE? $IPU�S�RETRAT��$SETHO�ST�en�DN�SS* 8�D��FACE_NU�M? $DBG_�LEVEL�OM�_NAM� ! � �FT� =@� LOG_8	,�CMO>$DN�LD_FILTE�R�SUBDIR'CAPC����8 .. 4� H{ADDRTYP�=H NGTH����z +LSq� D $ROB�OTIG �PEEyR�� MASK��MRU~OMGDsEV�gRCM+� 7$ �/�QSIZ�T�IMR� TATU�S_/!?MAIL�SERV $P�LAN� <$L�IN<$CLU���<$TO�P7$CCw&FRw&Y�JECZ!8%EN�B � ALAR!B�TP,�#,�V8 S��$VA5R�)M�ON�&��޶&APPL�&PAp� �%��'POR��7#_�!�"ALER�Tw&G2URL �}83ATTAC��_0ERR_THRO33USt9&!u8�� CH- A%�4MA�X?WS_Z1���1MOD��1IF� $�2M (�1�PWD  } LAطr0�ND�1TR=Y�6DELAC�0<%'�1ERSI��1v/'RO ICLK=HqM� /'� XML+ ��#SGFRM33T� /!OU33PIN3G_�COP�!�F�3�A/'DUMMY�1�G2?��RD�M*  $DI�S�SMC l5�M!n"%/7�ICC�%� FV�Re0GUP� _DL�VSPAR��S)N
#	3 _)R�/!_WI�CTZ_�INDE�3�POFYF� ~UR�YD���Sk  
 �t 8!]PMON� cD�bHOU3#EAf.af.a%f�LOCA� A#$�N10H_HE����@I�/ 3 �$ARP&&�_IPF�W_ O�F�PQFAQD0��VHO_� INF�OncEL� P����0WO�R�1$ACCEF� LV5[02��ICE�'p���$��c  ����Fq��
��
;p&PS��ADw# �5�WqIX0ALCUqX' dx
���F�����op�r�u�$.� 2�{ "���Qr�}�p�� �}��!�Mq5����$� _F�LTR  cy�p� ���������I�$�}2I��bS�HyPD 1�y�  P1�珴t ֏��7���[��� B���f���ٟ������ !��E��i�,�>��� b�ï��篪��ί� A��e�(���L���p� ���ҿ�ʿ+��O� �[�6τϩ�l��ϐ� �ϴ����9����o� 2ߓ�V߷�z��ߞ߰� ���5���Y��}�@� v��������M�z �_L3A1b�x!1.6�0���5��1F���255.�~�=���ܼu4�2 ;�M���a�s�������3��M�* ��������4+M�� Qcu���5�M�������6M��A�Sew���$RC��`G MA�� MA���Ѐ�v� Q�	 ���<-/b/t/G/��/�/�/�/�/�/��P �/"?4?F??j?|?�?@�?_?�?�?�?��? ��u2OLO�?wO�O��O�O��}iRC�onnect: �irc�D//alerts�O�O__ *_�EqOV_h_z_�_�_��_���sP�"��d���_�_�_o!o3o EoWoio{o�o�o�o�o"��$E_�o��(�o@iO:L^p��
��(�$"�r&J�u��q��� DM����$SM���ŋ��%1�D�� �I���8�q�\��� L�qN�q
!	�~������p������ #��USTOM' 
�}���# � ���TCPIP�r�}$H%�TEL��u !� �H!T�R�����rj3_tp�d�� (�ׁ!KCL����׏��v!CRT���W��"ߔ!CON�SX���ősmo	n]�ߔ