��   m�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����DMR_GRP�_T  � �$MA��R_D�ONE  $�OT_MINUS�   	GPyLN8COUNP �T REF>wP�OOtlTpB�CKLSH_SI�GoSEACHMsST>pSPC�
��MOVB RAD�APT_INERzP �FRIC�
_COL_P M�
�GRAV��� HsIS��DSP?��HIFT_ER[RO�  �NA�pMCHY SwARM_PARA#w d7ANGC �M2pCLDE|�CALIB� �DB$GEARz�2� RING��<$1_8k����FMS*t� *v M_LIF ��u,(8*��M(oDSTB0+_0>*�_���*#z&+C�L_TIM�PCgCOMi�FBk yM� �MAL_��EC�S�P!�Q%XO $PS� �TI���%�"}r $DTY?qR. l*1END14x�$1�ACT1#4�V22\93\94\95z\96\6_OVR\6� GA[7�2h7�2u7��2�7�2�7�2�8FR�MZ\6DE�DX�\6CURL� HSZ27Fh1DGu1DG�1`DG�1DG�1DCNA!1?( �PL� �+ ��STA>23TRQ_M���/@K"�FSX�JY��JZ�II�JI�JI��D �$U1SS ? ���6Q�����+PVERS�I� 4W � ��GQIRT�UAL3_EQ' 1� TX  
��(P���_�_�_ �_o�_%oo"o[oFo�ojjAQ�o�m�,'� k�� o'�������B�-�_�o�o�o�l�/VSe�k ��r��������d�#�5�G���=L3��R�y�?�z���@�����я���� �+�=�O�a�s���� rU������ޟ:T  2��!�3�E��W�i�{���������< ��ۯ����#�5�G��Y�k�}�������sP���$$ 1�\=�qE�� ῍�x���@��1�����Z��Wϐ�{� ��'�9ϛ����.�`�R�=�v߈� ���ߓ�t��������[sr[t>Tq� 6���Z�l�~�=�O�� �������� �2��� V�h�z�9�K������� ����
.��Rd v5G����� *�N`r1 C�����// &/�J/\/n/-/?/�/ �/�/�/�/�/?"?�� �/J?\?n?�/�?�?�? �?�?�?�?O"O�?FO XOjO)O�O�O�O�O�O �O�O__�OB_T_f_���,($1234?567890�_�U ���_�_�_�_�_�_o o;o+oGoOoao�o�o �o�o�o�o�o�o I9U]y��� ����!��-�5� G�{�k�������ՏŅ��$PLCLų��� Dm�?���1�%� T�m�x�c��������� �������>�P�