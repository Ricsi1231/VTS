��   ��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����PASSNAM�E_T   0� $+ �$'WORD  �? LEVEL � $TI- OU�TT  &F/�� $SET�UPJPROGR�AMJINSTA�LLJY  ?$CURR_O��USER�NUM��STPS_LOkG_P N��$�eT�N�  6 �COUNT_DO�WN�$ENB�_PCMPWD �� DV�IN�!$C� CR=E�PARM:� =T:DIAG:)|�LVCHK!>FULLM0��YXT�CNTD��MENU�A�UTO,�FG_wDSP�RLS�uU�@&ENC/�  CR�YPTE  ����$$CL(  ? ���;!��h D 0 V� IO� �:&+ ��>L!IRTUA� :/��$DCS_CO�D@���?%� � W�'_S  Jv*�!x �&�Ar91�"w!� 
 $B!���-�/ ? ?6?D?Z?h?~?�? �?�?�?�?�?�?OO�2O,#'SUP� `�+4OFO�#FfO�xO�O��  ��L�A���O � ��� V�[t&�+�j���D�ON_ ��W
_��+!�Ux_UCLUGH 1w)_ + �) �_�_�_oo)o;oMo _oqo�o�o�o�'�_�o �o�o/ASe w����o��� ��+�=�O�a�s��� ������ߏ��� '�9�K�]�o������� ��Ə۟����#�5� G�Y�k�}������� ¯�����1�C�U� g�y���������Я� ��	��-�?�Q�c�u� �ϙϫϽ�̿����� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������%