��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����DRYRUN_�T  4 �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	RESUME�_TYPENDIST_DIFFA $ORN41� 8d =R���&J�_  4 u$(F3IDX��_ICIDU�MIX_BG-yy
_NAMc �MODc_US�d�IFY_TI��  �MKR�-  $L{INc   "_SIZ��� ��. X $USE_FLC 3!p�:&iF*SIMA�7#QC#QBn'SC�AN�AX�+IN��*I��_COUN�rRO( ��!_TMR_VA�g#h>�ia �'�` ����1�+W[AR�$�H�!��#N3CH�P�E�$O�!PR�'I�oq6�$$CLA?SS  f�1���5��5�0VER�S��7 � �ץ1IRT�U� �?�0'/ �5�5��������0Ff�1E���%�19O��5OnO��X���5I2�;! �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_0�_�O+ W?�8�0 ��j�0*o�<oNi�� � 2~�9  4%�_�o��AA�o�o�o �o�o%7[��@�AM�=���8����dcs�yjc�$"+ uk"K�0��U�A`�XA�1�0 $N��������Џ�� ��*�<�N�`���F Au�A������ʟܟ � ��$�6�H�Z�l��~��4MbjcC!2ulu�ۯ���� #�5�G�Y�k�}����� ��t�ͯ���
��.� @�R�d�vψϚϬϾ� ɿ������*�<�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� �����,> Pbt����� ���/(/:/L/^/ p/�/�/�/�/�/�/�/ rv