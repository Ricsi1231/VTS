��   v1�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����UI_CONF�IG_T  � E$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]5�ODE�
6CWFOCA �7C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_Gv!k FKE�E ��8C�&USTO}M0 t @;AR$@PIDDbB�ChD*PAG� ?�^DEVICEބISCREuEF���}GN�@$FwLAG�@  &��1  h 	$�PWD_ACCES� =EFB�S�:1�%)$LABE�� $Tz j��@�32R�	�CUS�RVI 1  < `'R*'R�(Q7PRI�m� t1ކPTRIP�"m��$$CLA�@ O����Q��R��R�P\ SI��W�  ���QIRTs1�_�P'�2 L17�L1A��R	� ,��d?���a�P$b�da��c��`?�  ����
 ���Q�o�o�o�o�o�o�o �o( :L^p�o��� ���}�$�6�H� Z�l�~������Ə؏ ����� �2�D�V�h� z�	�����ԟ��� 
���.�@�R�d�v��� �����Я������ *�<�N�`�r�����`TPTX���&���˿` s�����$/sof�tpart/ge�nlink?he�lp=/md/t�pmenu.dg ��2�D�V�h�!��Ϟ� ��������u�
��.� @�R�d���uߚ߬߾� �����߃��*�<�N�X`�r�����Q[fq=bOb�� ($���������������Qa:�<cI�<gb�$�Bk
��\a��>ae����  ��\JP���������`�[`^�W`  �x�� ��S�QB 1�XR �\��_?b �REG VE�D��FXwho�lemod.ht}ml	singl}�doub��trip�brows�t�Y� �CUgy��C-gydev�.s�l/� 1,	t0/�/�� /�/�/m/�/�/�/�/?8?� �PP?b? t?�?�?�?�?�?�?�? �6�@M?"O4OOXOjO |OKE;	3?-?�O�O�O �O�O	__-_?_Q_c_ u_�_�_�_�_�_�_�_ �oo3oEoWoio{o �o�o�o�o�o�o�o /ASewE?� ������0�B� T�OOx���Y�k���ҏ �O�O���'�9�b� ]�o���������ɟ� ����:�5�G�og� a�������ůׯ��� ��1�C�U�g�y��� ������ӿ�� �2� D�V�h�zόϞϰϫ� ���ϵ����.���� ݿv�q߃ߕ߾߹��� �����%�N�I�[� m����q������ ���!�3�E�W�i�{� �������������� /��j|��� �����0B #x�A�S�9� ���//'/9/b/ ]/o/�/�/�/�/�/�/ �/�/��??G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O Y�O�O�O�O_ _2_ D_V_h_c�_�_m__��_�_�Z�$UI_�TOPMENU �1�Pa?R 
da�A�)*defau�lt�O�M*level0 *�K�	 Ho60�o�/o�o�btpio[�23]-8tpst[1�h�o�o�oko�}o(=h58E01_l.png<~/6menu5^yUp�q13^zr]z}t14�{l)q���� 
��.�@�R��B�{��������ÏՏd�p�rim=�qpag�e,1422,1 ܏�'�9�K�]�h���@������ɟ۟j���class,5�@�+�=�O�a�l���13h�����¯ԯ�m���53�"�4�PF�X�j�m���8� ����ɿۿ�l��#� 5�G�Y�kϖI`a .o��Rm��+q�������fty�m�o�amf�[0�o��	�c[g164�gf�59�h +q�ߣ�yx2��} �ҙz��w]{��s�� ��n�������� �����"�4���X�j�@|�������A���2�� ��/A���w ����N`�� @$6H��	�1\�@�����M���?ainedi��/�/)/;/M/H�co�nfig=sin�gle&��wintp��X/�/�/�/�/ �Ja���/?Se?% ��E?W?i?|?�?�?�? �?1?�?�?OO/OAO SOeOwO��O�O�O�O �O__M�>_P_b_t_ �_�_'_�_�_�_�_o o�_(oLo^opo�o�o �o5o�o�o�o $ �oHZl~��1 ����� �2�� V�h�z�������?�ԏ@���
��.��N�� d��������ϑO��5�As�̟�'�ٗu� ���� �����3��ڂ�h����̩6ٯu7� F�X�1�C�U�g�y�ď ������ӿ�����π-�?�Q�c�uχ�f"\1k��������	� �-�?�Q�c�u߇�� �߽���������Z �M�_�q���$�6�6����������d$�74$�U�g�y�������,C���5	TP?TX[2096��4��246�������186 "�B��
0�25��1��U���tvԡ���� i2�0*11����C:l$treeOviewy#�3C�&dual=o�81,26,4 �����////A/ S/e/��/�/�/�/�/d�/&�;x�53� �E�O?a?s?~/�?�?��?�?�?�?�/?�2'?�2��WOiO{O
O4�1%?>E���O�O�O� �6�O.�edit��O�OT_f_x_'� w5�1_@C�_�_�_o ��o4o�<o�Uo {o�o�o�o�o�o�o go/ASew� �������"� 4�F��?j�|������� ďS������0�B� яT�x���������ҟ a�����,�>�P�ߟ t���������ί]�� ��(�:�L�^��� ������ʿܿk� �� $�6�H�Z�	oo��?o ���������� � 1�C�U���aߋߝ߰� ��������	��@�R� d�v���������� ����*���N�`�r� ������7������� &8��\n�� ��E���" 4�Xj|��� �S��//0/B/ �f/x/�/�/�/�/o� ���/��?���=?O? a?s?�?�?�?�?)?�? �?OO(O9OKO]OoO 1�O�O�O�O�O __ ]/6_H_Z_l_~_�__ �_�_�_�_�_o�_2o DoVohozo�o�o-o�o �o�o�o
�o@R dv��)��� ���*��N�`�r� ������7�̏ޏ��� �&��/�/\�?���? �O����ǟٟ���� !���-�W�i�{����� ��ïկ�O��0�B� T�f���x�������ҿ ������,�>�P�b� t�ϘϪϼ������� ���(�:�L�^�p߂� ߦ߸������� �� $�6�H�Z�l�~��� �������������2��D�V�h�z���:�H��*default���j�*level8�M��	��� tpst[�1]	KyPt?pio[23R6�HuP�����menu7_l.�png��13��	5
��41u6�
�w�� �����//+/ =/O/�s/�/�/�/�/��/�/n"prim�=�page,74,1�/?-???Q?�c?n"�&class,13h?�?�?�?�?�?u?�25�?"O4OFOXOjOm#|<O�O��O�O�O�O�/218 ?)_;_M___q_|O�26x_�_�_�_�_�_���$UI_USE�RVIEW 1�J�J�R 
���_v�0oBo�m`o�o�o�o�o �oto�o+=�o as���To�� �L�'�9�K�]� � ��������ɏۏ~��� �#�5�G��T�f�x� ꏳ�şן������ 1�C�U�g�
������� ��ӯ~�����v�(� Q�c�u�����<���Ͽ ��Ϩ�)�;�M�_� q��~ϐϢ������ ��%���I�[�m�� �ߣ�F���������� ���.�@��{��� ����f�������/� ��S�e�w�����F�P� ����>���+=O a�����p �'9��FX j������� /#/5/G/Y/k//�/ �/�/�/�/��/�/? z/C?U?g?y?�?.?�? �?�?�?�?�?O-O?O QOcO?O�O�OO�O �O�O__)_�OM___ q_�_�_8_�_�_�_�_ o�X