��   ?Q�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����MN_MCR_�TABLE  � � $MAC�RO_NAME �%$PROG�@EPT_IND�EX  $O�PEN_IDaA�SSIGN_TY�PD  qk$�MON_NO}PREV_SUBy �a $USER_�WORK���_L� MS�*RTN�   &SO�P_T  �� $�EMGO���RESET��MOT|�HOQLl��12��STAR PDIU8G9GAGBG�C�TPDS�R�EL�&U� 9�� �EST����SFSP�C����C�C�N	B��S)*$8*$U3%)4%)5%)6%)� ''S�PNST�Rz�"D�  �$�$CLr   �����!������ VERSION��(  ����!IRTUA�L�/�!;LDUI_MT  ��� ����4MAXDSRI� ��5
4�.1 �%� � d%O�pen hands 1����% ?:�? �"  13~�0Closeo?Ђ?�?	O�9�7Relax�?�?GOmO�9	�6j82oOPO�OtO�3�?�O�O&_�O�6� +O__�_;_�4 �F�_�_�_�_�[�3�� (@�_6o�_Zo	oo�o ?o�o�ouo�o�o�o  �o�oVS�;M �q����.�� R�����7���[�m� ���ߏ�ǏُN��� r�!�3�m���i�ޟ�� ���ß8�J���3��� /���S�e�گ��ׯ� ��ѯF���j��+��� ����ֿ����ϻ�0� ߿�+�x�cϜ�K�]� �ρ��ϥϷ���>��� b��#ߘ�G߼���}� ����(�����^�� [��C�U���y���� ��$�6�!�Z�	���� ?���c�u�������  ����Vz);u �q����@ R;�7�[m ���/��N/� r/!/3/�/�/�/�/�/ �/?�/8?�/�/3?�? k?�?S?e?�?�?�?�? �?�?FO�?jOO+O�O OO�O�O�O�O_�O0_ �O�Of__c_�_K_]_ �_�_�_�_�_,o>o)o boo#o�oGo�oko}o �o�o(�o�o^ �1C}�y�� �$��H�Z�	�C��� ?���c�u�ꏙ�� � Ϗ�V��z�)�;��� ��柕����˟@� ��;���s���[�m� ⯑����ǯ�N��� r�!�3���W�̿޿�� ǿ�ÿ8����n�� kϤ�S�e��ω��ϭ� ��4�F�1�j��+ߠ� O���s߅߿����0� ����f���9�K�� �������,���P� b��K���G���k�}� ������(����^ �1C����� �$�H�	C� {�cu��/� �	/V//z/)/;/�/ _/�/�/�/�/?�/@? �/?v?%?s?�?[?m? �?�?O�?�?<ONO9O rO!O3O�OWO�O{O�O �O_�O8_�O�On__ �_A_S_�_�_�_�_�_ �_4o�_XojooSo�o Oo�oso�o�o�o�o0 �o�of�9K� �����,��P� ��K�������k�}� 򏡏�ŏ׏�^�� ��1�C���g�ܟ� ן$�ӟH���	�~�-� {���c�u�ꯙ���� ϯD�V�A�z�)�;��� _�Կ����Ͽ��@� ��v�%Ϛ�I�[ϕ� �ϑ�ߵ���<���`��r�!�[�
Send? Events�S��SENDEVN�T��Q�u�� {%	��Data�ߞ��DATA���o���%��SysV�ar;��SYSV�w���wO�%Geyt�x�GET+����x��%Req�uest Men���;���REQMENU?���y�]ߞ� Y���}�+�����. ��d�7I� m����*�N �����i{ ��/��/\/G/ �///A/�/e/�/�/�/ �/"?�/F?�/?|?+? �?�?a?�?�?�?O�? �?BO�??OxO'O9O�O ]O�O�O�O___>_ �O�Ot_#_�_G_Y_�_ �_�_o�_�_:o�_^o ooYo�oUo�oyo�o  �o$6�ol �?Q�u��� �2��V������� ��q��������ˏ ݏ�d�O���7�I��� m�⟑���ݟ*�ٟN� �����3�����i��� 𯟯�ïկJ���G� ��/�A���e�ڿ���� �"��F����|�+� ��O�aϛ�����߻� ��B���f��'�a߮��]��߁ߓ��$MACRO_MAXX��������Ж�SOPEN�BL ���2��ݐѐ�_���~"�PDIMSK�f2�<�w�SU�����TPDSBEX�  K��U)� 2�����-�