��  N��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A-  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  RO�T�AIO_CN�V� l� RA�C�LO�MOD�_TYP@FIR��HAL�>#INw_OU�FAC� �gINTERCEmPfBI�IZ@�ME�ALRM_�RECO"  �� ALM�"ENB����&ON�!� M�DG/ 0 $DEBUG1A(�"d�$3AO� ."���!_IF� �P $ENABEL@C#� P dC#5U5K�!MA�B 4�"�
� OG�f �d�PCOUP�LE,   $�!PP_D0CES	0�!e81�!��R1> �Q� � $�SOFT�T_I�Dq2TOTAL_�EQ� $�0�0N�O�2U SPI_I�NDE]�5Xq2S�CREEN_NA�M� e2SIG�N�0e?w;�0PK�_FI0	$�THKY#GPAN�E�4 � DUMMY1dJD�!UE�4RA!RG1R�� � $TIT1d ��� �Dd�DP� �Di@�D5�F6�FU7�F8�F9�G0�G��GPA�E�GhA�E�G1P�G �F�G1�G2�B~�1SBN_CF�!O	 8� !J� �; 
2L A_CMN�T�$FLAG9S]�CHE"� �� ELLSETU�P 
� $HoOME_ PR<0�%�SMACRO��RREPR�XD0D�+�0��R{�T�U�TOB U��0 9DEV�IC�CTI�0� � �013�`B�Se#�VAL�#ISP_�UNI�U`_DOxDf7{iFR_F�0�K%D13��1c�C�_WAqda�jOF�F_U0N�DEL��hLF0EaA�a7bc??a�`$C?��P�A#E�C#sATB<�d��MO� �cOE � [M�c���dqREV�B3ILxw!XI� Wr�R  � O�D�P�q$NOdPM�]p�0�q�r/�"�w� �u�q��r�0DfT p =E RD_E�pIq�$FSSB�&$�CHKBD_SE�deAG� GD@ � "_��2C�� V�t:5��3� a_�EDu � � )C2��PS�`�4�%$l �d$OP��0�2�a�p_OKv�USZ1P_C� ુd��U �PLACI�!�Q�:�� xa�COMM� �0$D���0�`��KO]B�
`BIGALLOW� (KD2�2�0VARg�d!�1>B ��BL�0S � ,K|a��P9S�`�0M_O]�����CCG�`N��! �� ��_1I΀7`��$�� �B�p�1S� �CC'BDD�!�I
�7���@�84_ CCSC9H�0_OOLF��P��qMMF�ݑCHs$GMEAdP�d`T�P�!�TRQ�a}��sCN�~�FS3�p|��!/0_FB�( ��؄pG��0CFfT �X0GRV0��MCqNFLI�0UIRE�+��!� OSWIT=$��N�P]S�"CF_�G�� �A0WARNAM�`�!1%�wPL��Z�NST� CORx-��8`FLTRV�/TRAT TX�� $ACC7a��� |��r$ORI��.&�RT�P_SF~g���CHG@I��rTꠢ1�I��T�
`%��>� � �#�Q���HD��a5�2B
BJ; CL�F�3G�4G�5G�6G� I�e8G�9�!��COfS <� �����3�ŐOLLEC���"MULTI@�b
2T�A
1ҠO�0�T_�R  4� STY2�Rf�=r�)2f��7�#Ӫ� |A06$��``��ph��P�* :�T�O���E��EXT�����Ɂ
B�уQ �2 
!��a0|كR.'+�b%��� �"��/%�Q���6�d�qc��$�3� 1�}؍1��ɂM�� ��� !Ջ-� L0?�� 6��`=A�$JOBt�B�����TRIG-�  d�������6�-'`V��%��e�_M�.b! t�F� 
C3NG&AiBA� � ��S���/1���pD@�q��0��Pa`����<�"I���6tB$4��
2J��_R��gEC>J��C^Jq�D/5C~	N�����0�y �RfT#� !������bG����HANC��$LG t�|�da���1��!A�`��xzRܱ1`��#�p>$$DB�f#RA�#AZ�0�jELT�� �PFCT����0�P��SM� �I��1� D��D��␶t�$����/0S��E��%�MaP
B aǰ�#HK��AE�0�����Ҡ��$  I| �sa�CSXC<���!% x�q�3��T�$_ПPANN�,�Y�MG_HEIsGHc��!WIDh�AVT�0�\�F�_ASP����`E�XP�1���%�CU+ST�U��&�E5b�%#IOv�-��BG_�`�a��' 1\ࠗ!�`OR�cK2D`ms���PORBِ �`� �aq5�`���P�p����0Kq11PXWO�RK��(Ϡ$S�KP_�`b�ѠDB�BqTR	p ) �! �P�ЬӰ�~�3 3DJ'dN�_CT��R�3��7PL�S a�dD����DQA'G]A�"�F����@@�`p &R DBt��*�231PRf�=�
�0�Q����+ ap��$nP�$Z��L�I!,�O�Cݰ��-�O�DeC��.�Ox ���9E���� /�OS�i@REs��B0Hz� C{R+$LKS�,$�C�^\[IN�EF�j1_D�j�RO�`�����������R���0�VPAɃ9uR�ETURN�Rd�MeR�U4�{�CRzP�EWM,0�SIGN��A�"!4qe��-$P�.3$P�Q�/`=�!&`:dQ�>`D{`R���uTaQ<bF�GO_AW���Pp+0
�&!��DCS�pm�CY-�1��`1[��a��*�d2�j2�fNQ���x�)�cDEVI�P� 2 P $fǶRBE���PI�gyP��vI_BY���&p5wTJA�dHND�G�A3��jcsE8��d�� SBL'�˳Ђs�d�A�bL�4� Hf�y0���fTO3FB�|%�FE�Q���r�d�cv&5�rDO8!V�=�MC��]�F Pz3'��rq�H�Wߒx�3R�aSLAVQ;6��INP��5v���k��ao�7D *$DIS� 0\�0!�0��Ơ�������̃�:1��:1W�P�̂NTV�ӧ�V�ð��SKI�TE�`v"��%�Z�8!J_�"_�@O�SAF�E�`�_SV��EOXCLU��a0pDi0LP���ڐv"�֜�!>�I_V�r�P�PLY@u���DE�����_MLQ�a0?$VRFY_�3��M��IOt ����P��Z�Op��LS(�P1"YD42�<��c	���0P�5k��`�AU��NF/&���ee��`Q�#Dw�pM��Si���AFK�CPpP���q 8PƲ0TA�0�� ��t_SGN��9 I����Pa�#���!�>`�1��2)�� UN��@��Q��e��'a0 `	 q�n��v���/2�EFv0I�B: @b�pFS�4��OT` _�YD1AYD?AG�VA�0[EM'pNI�B;��� �A���DA=YP3LOADtND���ZC5VA�EFV� XI�r<PDA�3#O^�S�0_RT;RQ��= D�p<P���Q_0 ��E�`��^ŭ�< �a��<��_��AMP� � ��>:��¬�����Wc���DU`����2C�AB��?��PNSl����IDh�WR��h��:�VwV_��~��> �DI�����@� /$V`SEQ�T5��N�ypO���1@��BE_l:���VE���SW�щ�O -С��2��=� ��OH����3PP����IR,1��B�0<��Ã�
b����)�BAS��$��w#�vխ�?����p�ތ�RQDW�MS�>���AX�׳���LIFE�0����`A��N������n�����Ch ]�n�C& aaNA��!t�n�OV����HE���SUP$k�@����0_;��B��_��]�zai�Zf�Wf�&!i��n�sr�cXZCA��Y2��EClPT�0�P��N������� X$A `�pM HE7SI�Z�� �bN�U7FFIe����0�L�NDW�ZC6��fAM�SW��B 8z�K�EYIMAG�STMmQ:��Q�i��!����VIE��@QC ��uL��ÃC?���� D��mA�STO�!� 1@�?@�L��W�� EMAIL��P'��hн�FAUL�BEp��S�3� COU��� ��T:P��F<' $f�S��9�;IT�sBUF ÁP �d00:�B�� tC��g,3tSAV����������s0r�P��=P��p_���9)OT�Rg���P��G@]*��`'AXP3�!� �_��#_G��AYN_�APG��DuN@'uU�M��TW�=F�P�E�0:P$�@QHd�9&�wQ��!���p�R@QI�0GP#1ZA#C_�P�PAK�TE0*�@4\�R�8?5K#1DSP�#2PC�;IM�}3�1ĥ#1|�UZ70�U��>IP�#3�D  |4TH7@�sp2c�yT�Q}3HSDIz6�ABSC���PV���-J+@�#3DQ`s�NVv�G\C3D��z6�	F�Ѫ d_3� �!�Q�SCn�u53MER|��#1FBCMP���"0ET��APJyFUN�DU���`����CDs9�0T O!0OR_NO��@QK����`R�T?�PS*UC�0+UCh��!��!Sg 
�LH ��rR��rS�F��h� 2��TBa�VVL��VPW��Vc�V7�Y8�Y�9�Z���X�Z1�Z1��Z1�Z1�Z1�Z1��Z1 j1j2j2T�[�Z2�Z2�Z2�ZU2�Z2�Z2 j2j�3j3�Z3�[�Z3��Z3�Z3�Z3�Z3� j3j4b�0�EsXT�	�M <(�  X� ��� �U� �w@U� 0FDRn�NTrVb�["��%�\+B��REM��F�QN��OVMV3K�AT�oTROVT�DT�6t�MX��INT��s�k�IND����
x��@� $DG�! 0�}�� ���D��}��RIV�@����GE[ARV1IO��KD���N� 2�^��譐� |V���Z_MCM��n���F1�UR�B�O ,)Q�?� �0?����?��E����Q���@�P��s�Pz!�{�RIU� �ET�UP2_ Q L��TD�07��5�਑�����q�BAC��"R T��	4)�:%��aS� �@IF�I�� �@�P��P�P�T0" �LUI��S � �	hUR@���?2�!+@�T�Ө�I8�$̢S���?xؠJ0CO�, O#VRT�p˰x�$SHO��}�PASS@Z!���0���jG�Af�TFFU{�	1�!A�22����f�wU |΀NAVj �̠�u���><��J�VISI��I�SCr��E���Ѫ�V��O>�o�B���E�¶$PO���I��F�MR2�V $�P2�%�0�)��0�B�T�k�V��D�_a����_z��D���M�� �DGCL�F�DGDY��L	D���5�����ڑ�M`�W0[�� T�FS7 �X� P�p7�3� $GEX_7�N�7�1� �y@�8�3p�5p��)GGA�Y��
����W�Oy�DEBU1GAs��I�GR�(0�U�CBKU�@O1nn` ��PO?�������@����M�L�OOz#�SMk�E��+�����_E �Z � �TER�M@�[I��ORI��!E�\I�`�SM_0�E�]I�3�6����^b��@UP�_�� -����Z(̠W���[��G�����ELTO0$U�SE�@NFI����{��є n���\$wUFR=�$P0��2��Ev�OT?�b@�TA@%�Q�NST�� PATA g�P'THJ�A�@E� "�@��ART �V8!0��REL���!SHFT�2��m��E_�R�@�C�� ��	$����^��&����3N�"SHI���U�R= �AYLO�0�! �!�����m�b�3U�0ERV�P8¢���r M�� ��Aql���Ql��RC��3UASYM�!3U��WJ��qĀAEȓ���	¢�AU�@� �!��V�E��P�3XU fAOR� M ���/��`=����0l�,�!�HO�ԇa �S�p�۰PO�C����a�$�OPg����)�bR�@���@��R�zC�!OU-Cm�e���Rk�����<�eo$PWR�IM�iR_�����������UDȒ�p��$b��$H5!z AWDDR�vH2�Go�(�!�!�!TPR���c H�pS�@��As��%�S�%�S�%�SSE8+Ѱ�7��HS�@��d $?��_D��p���2PRM_�r�SHTTP_�PH�e (�@OcBJ���"<�$�v�LE^�:4@�f �s �w�1AB_���T%�2Sy-C��K�RL0)HITCOU,DB�L����2��Ȧ
��n��SS�À�TJQUERYO_FLA�0Wa���g� S@P	U����O>F�1�TUB��$VA�$VA�R �IWOLN,�h�@w��C�!$SL�$INPUT_��$��HP�FPT�@SLA�� i�@�O�E�D��E��1IO0F_AS:�j2�$LG�c7G���PU�����0�C�ЛC: HY�w\Q�5SSPUOP�k `!PzQ�v��LT��SV�Q PF#��W�Q�SV�R�Vr1UJ�lo �  �NE��+��RD�D�J7z0O$J8&i�7p�I�/bAg7_LAB_�1`Yh%aoAPHI��Q0c:ugD9�J7J�q�p�^�_KEYʀ ��KW@LMONz�m�p$XRP�K@�sWATCH_pΐRF��QELDI�gy��c�n ���U�V^ �v
rCTR`��
rA���@LG��o� !�yLGŠZ���Wu�VvPVvFDaxIUxlx� cvTxB�VvSp��!� ��P��p�B����������_m�E��`�&�[�Fa-�G�Spr�(Rq^q�l��l�Pl��px�I�k�����l�B�l�SpRyS�`|�  (��SLNa�p�P�0@��`��B�`�q�U$3���yL���DAU�EA,0W@�4�*��GH�r1$PBOO>,�q� C;R@ ITCh���7V��}��SCRT���<QDI26SS,���RG��� ���F/S�ݒ�4$Q���,VW��$Q�/SJG=M�MNCH!B#R�FN�b�K<�PR�G:�UFH���H�F�WDH�HL�STPH�VH�q�H�o�H��RS��H/d�,VC����/S���U #1\���� pDSO�G,���ݰ,V�������(�2�OC��K�EX.+WTUI:�I�p�ǲ��ҳ�ҳ8�<����A��	$����;NO˶ANA$R��Ε�VAIY`�4CL����DCS_HI��O��#N�OTȿ�WēSIy�k�Sw�ҘI�GNlp�@~s9�@TܼN�DEV�LLvaV�_BU�Ъ@�rp T��$bwEM'WGAt5r*��Ap"sp �@PQC30��n�1F�2F��3F�や�O���t ��P�8;��D���DIDX���Dn����Z��ST{PR5�Y�2p���� s$E��C�ۓ0"0���p1�h�P��u L8@ J_�_X��'W�!D%�EN,0D$fԚ�_ v g�20rB����� �MC��w ��PCLDP|{P�TRQLIj�p�	`���FLG����]��>�D�a��)@�LD������ORG 	`����gE��#g��"��]x � �	�������SwTD��`��.����RCLMC��I�[���{@���@M�0Q_��y�`$DEBUyG�%DATA�r�5T4��3UFEB`=T���MI� ]gz d����RQ�`=��DSTB� ��c sˑ�AX���`��EXCESH��VM ^�{0�g��j0U1_�|
6@u_/ q�P����K;t} \�8@'b�&$MB*BL�IS1aREQUI[RE��MOfOv�����L`�M�e~ 0<Q�1rT��ND
�Sp"���x�D7��IqNA0���RSM`(��N���q��S��PST�0 �nv"LOC��RI��v��EXt&ANG�Ҽq�ODAQ�e��c $�`���bMF F���%��_�K�i��%��[SUPe��F�Xk IGG{� � ���_��q��_��_��`^`%��'9{P 78{PF6'DS,�, EE�0E2qC�pM@n� t� MD�1I>�)�6���4��7qH� *a�4DIA]a�3ANSWᑽ4,�T���5D<�)��O�Sܡ�_�� � CUBlpV�0��qO�A9_ ^�� ��P�C��# �y�pnHP�nN +`u@PmHKE8��`a�-$B�PaF�QPND2���c�A2�_TXh�XTRAh���B����LO6�b_��� To �F��R�5B VS�RR}2�U�0 #Q��A�� d$C'ALIy �uGB�\W�2��RIN^�`S<;$RjPSW0���S���ABC�(D_Jp�@�q �1_J3�V
�R1SP(pD`q 	P�T�]3�]:A� q �eJ��%ej��O���IM���CSKAP��Td3��TdJ=���QTl�eke�e{g} �_AZ��!a�aELx�� b��OCMP�#������RTA�cUc1�"` U��1�xt�zZtSMGѠ�0��JG��SCL<� x%SPH_�����s�Xs�@cPgPRT�ER�P`S �I-NxpAC/҉5B�udՒqT�q2�_N^���u�r�ѫ�z�t�͋�yDI�a�q ��DH� �@^��5��$ViP#Qs�$@/p<�C�[Ќ��A���R(C_��H ��$BEL�`�uq__ACCEL��W�|��f�IRC_R�0���<�NT�ѳ��$PS�p��L   e�����p|���C�}� �A\�҇r�҇3��F0�_C�&��	���-��C��]�_MG̑�$DD&�}���$FWx�0b�B�r�]��7�DE`�PPABmN��ROYpEE� Gѐ���{aG�]�~��$USE_hPJ�P�@CP��Y���8��� 8�YNY A l`�D`�1�M6@A�� �OL�INCD�!_�F��?�Ka�ENCShP|1q���]�~��IN��I𡂆��0AtNTVEx$�`S��23_UVa��Ҵ�LOWL�� ���0��k�ԦD-�q [xpd�k�C�p��MOS��,M@	�����PERCH  �O�@{r 3��!>� ��ע�����g�bڕ��$��BcA����L�Bc�)Ag��� תҶ�T3RKyu��AYS�� ����Æ �fM���MOMB� ?�:@o^�\W�ԃ�F�7�DUJ`��S_�BCKLSH_C ����6 ��@��EB���f����}eCLAL�К�<C�� ��CH�K���S�RTY@b0�C���51�1_��N�_UM/B�C/p&�LqZӛ�LMT�P�_LC��cs��1~�E xݙЋ�wЎ��Վ��P05����w�PCD�w�!Hf��*�B�C���D\F�8�CN_wRN��L9���SFJ�h�Vڒ�)�|�uqᡂ}��CATI�SH�#wR8� n�1�}�}�U��Ypf'�PAI�=�_PH�,�_X`Lp	�'�Wa�+��JG��� � �OG,�p�TORQU̐�U�"�n�W�q�n���_W[��q@'���������I��I��I�F� ��,bX;a0�VC\�0zr$1*� >�1�JRKNob��D�BJpMfC��M	 _sDL���GRV��`�����H_S8�Հ�
COS��`�LNq Q� /p��J8��1Z��MY����A��THET=0ݥNK23��lQsCB�CBQsClPAS+!���!�!�SB�)"�'GTS�a��C�Q�!�w��w_*G$DUж��"\RI�1�&�Ka_�Ql2��_�NE�Zd� I*��i�w$�p�A��%�'���LPH��"���"SQE38E3G�"VPo3Y:v�pV8V8T�.<V=:VJ;VX;UVf;Vt;V�;V�9H8�65B-=��LHJ;UHX;Hf;Ht;H�;UH�9O<O8O�I�,>O=:OJ;OX;O�f;Ot;O�;OvF��"�TY8YT	7SPBALANCEd���LE@ H_�S�P�q)�R8�RGPFULC�X�R�W�R�G�z1��aUTOy_�?�T1T2iX�2N��c���8d?q@<��P� ��S�W�Tð�O�`e���INSE9Gc���REV]f��Ε�DIF쵾y1�l�g�r1���OB�a���i�2z�ї?LCHWAR��ߒ�AB��k�$ME�CH!��q*�AX�P��.v�'�r`�� 
/r���~�ROB'�CR��qu#�; 5�SK_�P;�_� P #`_ʐARX���t���1|‧����p���ģp�aI�N~a�MTCO�M_C ?�� � !��`x�$N'ORE��
���`�ro� 4f�GR���uFLA~a$XYZ_DA
1ǐ��/DEBUA� ���&�� �P$�COD�� q�@�p�;�$BUFI�NDX�� `�M{OR�s� H�p Y�g��Ƶ�7���ėb�L�(�Ɇ��T�A����`�i�G���� � $SIMUL)�x�Z�������OBJE�P�AD�JUS3�&�AY_�I@�|�DT�OUTpI�@�Y��_FI�=��T�������� K��`*������`�0���D�FRI��˕T&��ROi���E��ΰ��OPWOp �p��,~�SYSBU<�0��$SOP�������U��`PRUYN�r>�PA�pD=�r�u�_o���3��a�ABeq��o�IMA�G���p� P�aIḾ��IN� f���?RGOVRD��/���q�Ps���z�^`L�_`���>�Y�RB��з���MC_E�D��p ��N�@Mx��ш�MY19��7����SL�P�p�� �ZpOVSL�]fSDI�DEX B�T�Q�ñr�V��o�Ny���l���w�����'���C{�TJ�����<���_SET��p�� @f�ڲ8u��R!I���E��_!�����^��a1�n� 嗯�Tp>�ATU}S��$TRC� 8����M�BTMV�@�	I[�%�4��,���p� D�pEo�X�J��0E�bK�������K�EXEQ�+���¹�Ą�ⳙ鰡pP�UP�K���ɰIS��XN�Nv�Q�%�y�	��PG�u��$S�UB?�8u�?��J_MPWAI��P|��W�LO��;��`��$RCVFAIL#_C�q"�Z�R��"��+s�l�C�up�ՅR�_PL�DBTB8>�p�"�BWD���3UMn��IGV���>a��TNL�����ҁR���7�}�|�� P�EED��R�HADCOW>�s��E]��K�l�)�DEFSP>J` � L�p5p�h�_k�9�y�UNI�t�{�w���R��ƳLT��`PI�ֱP�p�q�m�g��s���L�t�PǢN�PKET�┛�Y���P�ҙq�� h s SIZAE��<���K��S1��OR�FORMAT`��CO7��b�EM't5���UX8������PLI�ҙq�� $�OMP_�SWI�`^�EB�W�"�#��s ����AL_ ���v�ۀR��B��C�rD[��$E���J3�D��� T�PD�CK��&qǢCO_J3+4��
}R�q��6��	���C_����� � �!`PA�Yw!�r`_1g
2g��J3t �s����TIA4�	5:�	6�rMOMƀ�������pBn�A�D���PU NR�.�.��a�z�t�` I$PI�&`�ql� l.#l##l$���"$t$]�R&l�R&��}q&w���/�HIG ��/�o�h�"&h�oե� ��"&X#1(��@)��o�SAM�P���$"'�#No�MOV���`�p �!�`��r�$l��&h� t �)� �r� �%d��H>`�#IN#< ��x#*8F;!4o�,:l8xC4l;�;GAMM�V|S�K�$GET�����=�DP�
3`L�IBR���IV�$HI��_��Y��rF�EۀHAN+@FLWMIF@L+ImFFL'v��C���`Π�o ��I_w  �脮�a��5�G����I�� ��$�� 1�o�I
�R$pD�c�b�����`LE�q�q�bXL�*P��MSWFL���M��SCR�7 n��V��U�Y�`�p7�PsaUR�W�Q�/��S_SAVEc_D��U��NOP C���Q�P�4`� h	��h	�hjXk�$��h�Db�v �2 ,��&�'�"�s(�,& ȡX(�g�e�c�!�����y�M�u� � F�CYL~��7сS����Kwj����SWs�����P-qW*`�r�rN�s�-qM���{CL�x�E�$(��X1�x�M�Q�?� � $Bq �$W�L�ʀ��� �(	�/	�6	�����ȃ�1�0������X��O7��Z��x�B�n�� ��AOMSj=oOoaoso�o� �CONURȠ�SP_/ҧ |��ň�P�	 U��U���P�
��m���
���5)�)r9��R��)�� 9�P��P�M��QU�  �{ 8��QCOUQn"�QTH��HODrn �HYS<�ES�!F��UE��R��O~��  ��P�p�5�SUNR�ws*pO"��� P��J����Q|���ROGRAe��Vr2��O��I�ITxXP��-�INFO��� ��}���Vr�v)qOI��� (�pSLEQ&�%�̀�c�OS�@,��{ 4��ENAB7�>��PTION�K�p�D�_��GCF%�ů�J�Ю�Q����0Ry�E�W��O�S_ED\Я�� I����K�!� A�E>@NUҷ̸AUyTaϵCOPY�!P���_�#`MAN������FPRUT� Z�Nk�OU����_RGADJ���3X_-p��$��u���u�Ws�Ps�pPu��/�e�D�EX��YCn7��a�NS!�9�9p�PLGO�C� �NYQ_FREQ�EWw0&�J�G�L�AXS��s��w0��CcRE�0��@IF����NA�!%D�_G6�TAT��p��7MAIL�"�a��dP�������a��ELE�M%�� �,�/�FEASI2��b�"` ]p����a��P�0�0I���D����ƐgS&$�AB����E��/ 9V��<�BAS��=���2FUM ^�`�$T�p�RMS_TR��UP�㇃L �"`��p���«��D��	�� 2�  R3t�@4��z�����p�P{qz��x\TDO�Uv�PTN]���PR�p&���GRID����BARS'T9Y3�_�OTO� �W� :�_`�!����G�O��"�� �s ����PORv����p��SRVd�),����DI`Ts �������4	5*	6	7	8��)q�F�2%��8�$VALUW��U��0�Y}F!��� .��a����f��XR�AN�S�v�R����aTOTAL�#F��PW��IO�REGGEN�
��X}�`^��Ǒ��TRc�E"�_S�Pc��AVs������\�E���S���bI���V_�Hp�DA惃�S�_Ya���S�PA�R�2� Q�IG_SE��m���_M��C_{�eR���*�`� �=#(SL)G�%��q��RՐ]p�t� � S�r��D�E��U�Q?�,�r T�E�� �� !�<�B�JQ&b��IL_M&�� eS���TQ��3��w�WzrV!;C/=P�0��93mMP9V1O:V1];U2l;2];3l;3];4l;4]:�Q��C�P����6�q�bIN�9V�IB�p)4@�aD2�H2%H3H3%H4BH4%H���S�R����D $MgC_F	��@�`�L�Q�Q��M(`I�C�B(� F�!�`KEEP_H/NADD�A!�DA��IC��d��D��B]p�COߑ�D4��A�`p�Cw���CREMR��D���9UPQUXU�`�e�DHPWD � �CSBMS�K��COLLAB��t� �P�J�ؠI�T��~���E��� �,�pFL4�a`Y�N�@�\M��C"�~ UP_DLY�=�8�DELA`�Zs�YƐAD����QSKIP0u� i���K�OY�NT�1{qF`P_K�t�eg|� s�$�|g��i���i  �j* �j7 �jD �jQ �j^ �j9���J2�R�����*�Xb�T  �+q���+q���B+q����AC`RDC��+ ��Rz�R�(0�AR9�uz�tr��R�GE���|s?�FL�G��|�����SPC�����UM_+p�#2/TH2N+��pp� 1�  ��S�11��� l`F���Q/��SAT2P Z�� G�
�E�����<� ����;�Q��qHY�f�W ��2���`.�@�R�d�v� \p
�3�ř�����Ϗ(���4���(�p:�L�^�p� �5�Ǔ�����ɟ۟V� �6���@"�4�F�X�j���7�ɍ�����ïկ�|�8��
��.�@�R��d��S�P���@���)�p�RPE���9 �p���IO�!<�IŰ� ��POWE�1� Q��PIq[qE�� ��Uw�$DSAB�_б��`C�p|�c RS232"�'� �mp��	P� �ICEUV�u�PE|��PARIT��u�OPB�P�FLOW�TR��aQ�8�CU��M��U�XTA�P�INTERFAC��x���SCH��� t`�@�@�� !�q$�&�OM��#A�p���I�Cm�
�A�#c�T������Xm`�؎�� EFA�@�B�Q�kG� $a_� *3�x A���� ��o�i  2� ��S`p��	� �$�p,e�r�=�r� _�H�DSPT��JOG��C _Pra"�ON p.eqp� z4�K��_MIRp�̐�R�MT3��AP@3R��p����qS�ب��qPG��BR�KHgѪ��P�da �^#�?�P�и=㞪�BSOCH�RPN�D�D�Y16�a�$SV"PDE_O�P $FSPD_OKVR�A$`�PD�&��OR����N� ���F��m�OVp�S!F�� ���F����� UFRA��TO��LCHb.e� OV~��Pm�W
`�Vm��Q�Q�|�#  �@�rTIN��!/$OFSn C���#WD��1��P���j�TR���/!_�FDdS��MB_C�P�B`�B� �Q����SVKъ���_,c��G���AM��B_h�X3_�M� -��!8�e T$SCAc�� D�j�HBK�ѩ�IOⴵ�X��PPA �����>X�e?DVC_DB�"� �ѕ���R��%a@(X%3&^ �s4p=��5�~�U�#b�7�CABTp�'z��&���
m��_1Щ�SUBCP	U��z�S�p"0dS���a�)�t�da$HW_C��Жa���&�a���@|@��$U�P!�00A�TTRI��(2z�C3YC�0w#CAT"��FLT�0�0Ƴ��Z#���qLP��CHKގP_SCT��F_�7F_<�20:FS8���2CHA�q�7p�1�"��2RSDa`��1�ӕ�X�_T0P@ ��EM۰RpEM�T�2�`|@�2�bc]CDIAG��R�AILAC��BM `p�A�RZ��aQ^&X'Q^%*#PR�S�P� d��AC���	^WFUNCcb<�'RIN�p�R$oA�DLу`S_M��j�SqpxS�qxCBL�`$X@TA9[51<X5XDA�QzX@S9ULD��r��SU�Q�A�STI�B�U8��f@$CE_RIYA�q��AF� P����SP �UT2�@C���"�OI0�D�F_L�����L�M�FA> HRD�YO��x RG�PH�	@����PAeMUL�SE1`���'c�P�$J��J�����F�AN_ALMLVܢ��aWRN�eHA�RD!���vP2$?SHADOW+ ���I��b"�`��!��_,, �&AUL�R�4.�?TO_SBRX�Js�a�Sz0��AksMPINF�p*1~t�QΉsREG���aDGĤP�sV�И�	�DA7L_N�FL5dB$M�P�0z�� z ����$Ʊ$Y
���$��)���� ���EG0�@=�r�5�ARO�8��Z�2c�D�fP��AX�EW�ROBT�REMDT�WR> �_���6�SY�o��S���WRI> H�� SAT��U�/���E1AذQ��C+qM�B ��d�5�CDOTOr�qذP ARYT�`>��AD$뢆�FI��~5�$LINK0a�GTH]���T_���dP�6d�X�YZ�Ґ�7��OF�Fl ]���y�.�O	BR��B�4!���@�FIC0��=У�j��Bl�_J���җ� j�� p� �8d����&@4�bl�C����D�U�O�9�ETURB�`X�S��L�yrXπrT�FL�� s#B��à���30d�z W1�ذKy�M�$Z�3�!�B�%�B�'��ORQ8Fa�S��!�B��O����t���8_�q��OVE��
�M[�u�	����������qѧ��A��0��AN�!`����Q����� �,"u�������2���2�ͳa�ER~�Q	B�BE> �Cp�A�f@ �U3BJ��Q~&�QAXA�ҁQD �! _���cA�ɍa�ɢ@�� .��ʝ��ʼ���e�������1����A`��A` ��A`��A`�A`�A` "�A`2�A`B�A`R�o��c�DEBU�#$��A�cgB���AB��G��Vt�" 
.�#�V��!b� c�b�Ab�.�b睑b� ��b�e�b眡�Tq��R\_��LAB��T�� �GROm0T��l]B_AAW�선� ��Pp�?�U�;�>qG�AND�� e�^!��h�>q�� ]�p����0CQ��`0��NT�`5��VELGA���A~���SERVE��N$�� $�@PA$! POsf0� �8�����#���  $,TREQvr
+��5 �9��R2�J�P|@_ �� l�@vERR ���Ir���N�TOQ��Ls�P��܂�3@G
%s��2*p4� ,hNh ��RA�? 2� d�s �A  ���$��FB#`��_Y�+OCrQ3� � �COUNT� � )FZN_wCFG4� 4� �vf2Tt�"-!�� � ��I �� �S�M�0�b�N  ����0�FA�P��V�X��+��
�~��z ��Pu"K H�EL�p��� 5� B_BASN�3RSR�v�@���S1�Qx 1�x 2��*3�*4�*5�*6ʛ*7�*8�k!ROaO�0� d���NL��w�ABy@y AC-K?�IN=T�0�r�$U px`�1+9_P�U�3�`�2OUP��@�xX#��0�T�PFWD_KAR���q� REW`P8Z��QPQUE�y3@ ����ݢ�`qI�`B��X#���C��v��SE�M^�Fl�s`A�S�TY:4SO	@4tD�IF1�@��1��!a_�TM�sMANRQ�wF��END��$�KEYSWITCaH�3�1YA�4HE���BEATMsPE�E�LE�Q'��HUҝ3FD�2S^DDO/_HOM�PO�.0EFl�PR鑪���G5C�@Oca� ��OV_MF�
p�PI�OCMr��7j����Y#HK#�� DH���w�Ur�2M=�x�4ɰ��FORC�s�WARSbKY#OM>F� � @���=pU�PD�1�V2��V3�V4h�zBOʮ0L�R���xUN�LOd0t9dED�#q  �SNP�X_AS�� 0��p�p�q$SI=Z�q$VAE��?MULTIP2��[a�PA�Q� � $s9Z`R��m��S�-�C� �fFRIF��=S�0�Y!T��`NFzDODBU π���esynRy n$�� x� SI��TEޣc���SGLUqTl�Ϡ&�ns�<��VpSTMTܡ�s�P1���BW��WtS�HOW�u���SV�b�_G�� e�$�PC�>b���FBZ�QP�xSP�0AE0��uMVD�p���� ��A00 ��!��P)��P)�`)�T`)�5'�6'�7'�U8'�9'�A'�B'�@�P)���*�
�)�F'��b��3�1@�1M�1�Z�1g�1t�1��1���1��1��1��1�1ω1܉1�2�&�23�2@�2M�2*Z�2g�2t�2��d�T����2��2��22ω2܉2�����P3�i���M�3Z�3g�U3t�3��3��3��U3��3��33ωU3܉3�4��43�U4@�4M�4Z�4g�U4t�4��4��4��U4��4��44ωU4܉4�5��53�U5@�5M�5Z�5g�U5t�5��5��5��U5��5��55ωU5܉5�6��63�U6@�6M�6Z�6g�U6t�6��6��6��U6��6��66ωU6܉6�7��73�U7@�7M�7Z�7g�U7t�7��7��7��U7��7��77ωe7܉7�bVP�@=U2� ; �࢐"
�qr���P�>�R�1CM �Mb# Rd K ��Q_V�R��S�P��MY�SL�   � � we-r��dlgPf�x�@(��rVALU��P0�6��a�F�ID�_LzC��HI��I~�R$FILE_w3����4$S* �S�A1� h � VE_BLCK��3��pq��D_CPU	x`	l`������_��@r2R �? � PWX0l`gLA�qS0�l}vRUN_FLG�k�v�@��k�vHq0�� |vF�TBC2�_� � .`B� �S`�1A�@&D4CTDC� �'��c5"TH4&P��\�R1:!ESERV!E'C}4C}3�r� �30R �X ;-$�LEN'C��4C�T0RA�0#L'OW_�31���M2�MO��BeSpC0IY0��)���,+DE<%qLACEWR�CCAc��@_MA]`;&u%K'u!GTCV|,�!K'T�A �*�%�*�r:#�q�%K#��qJV1�uM4�0JH�7�:%'1K%��2?@�p	�@19#G`JKS6VK'Ae1iQe1̞Z0J0z4i3JJvq3JJy3AALi3P�0q3�0�64�55Z�@N1�,�0�+y ��L _�q�@��� C�Fab� `��GRCOUo�qq|B�qN�C�c+@REQUI9RhPEBU�c�n6$T< 2�aA�KF�``�� \^�[APPRW@C�@~�
$OPEN�HOCLOSP�HSE��I:%
��f� �M7z � Eb�D_MG�QPC���X��P� WBRKYN�OLDV�pRTMCO_WWA]UJ`PSTP�4W q3W y3W �3W �3W 6�Ucq�R��p >qUA��G� TB���W<q1�SPATH�Wa@ca�c�`f@��p�qSCA�BWW�BQIN�UC ,qg`-C�UMphY��c vb���jq0�j��`�PAYLOAOWJ{2L��R_AN/�cLh �i�a�i�aUR_F2LSH8rtLO�dfaw�c%w>�cACRL_��de�Wp`g�dr2Hb���$HR�rFLEX�C�J�� P@�B|� E�q>�� :�� K �.��s1K ���F1.�|���// )/;/M/_/��Ei/{/ �/�/�/�/�/�/�/�� ���'3S4��Ƙ?,?H>?-�E:T����X� 1Q5��\5e�>�h? z?�?�0�5�5�5�5�?��?�?�:�rD� ��� O.O@OM��AT��SA0EL��{�jZHJf@�a@JE>PgCTR`a��TN���w�KGHAND_V]B��$�@AH�� ���P���  � �ٰVER�SION�������IRT�U�p���AAVM_WRK 2  �� ?0  �5�W�rc�Tφ� ��A	���ͽ��!�������������ߨ�`�S�e�m�1�BS��� 1�� <A߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZl~����8}�"�(�LMT������  d�I�N���PRE_EXE(3 &�`�n���� �1�IOC�NV�% ��P�[&US'%��|�IO�_`  1>�P $.�����-"ܻ/!�?����/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p�� ����� ��$� 6�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲�����LARMRECOV J%�"��$LMDG �'� �LM_IF �+��q� �����_����������, 
  �H����,n��������3�ANGTOL � J* 	 A�   �����PP�LICATIONg ?J%3 �3��Handl�ingTool �6 
V9.0�0P/03���?
88340:M
sF0s`5458�M
BT7DC3xH ��6None���FRA�� �6��P_AC�TIV�)�~UTOMODF �*�)P_CHG�APONLD �XOUPLED ;1�)� �����CUREQw 1�+  T���	/)% �>$�"��3*$H���#*HTTHKY 7/�+//�/�/�/�/ �/�/�/�/??/?A? S?e?�?�?�?�?�?�? �?�?OO+O=OOOaO �O�O�O�O�O�O�O�O __'_9_K_]_�_�_ �_�_�_�_�_�_�_o #o5oGoYo�o}o�o�o �o�o�o�o�o1 CU�y���� ���	��-�?�Q� ��u���������Ϗ� ���)�;�M���q� ��������˟ݟ�� �%�7�I���m���� ����ǯٯ����!� 3�E���i�{��������ÿտ����E#�T�O��$6DO_C�LEANe��N/M  ��5��������0��_DS�PDRYR��H	IB��@�Ϟ߰��� ������
��.�@�R�8d�v�MAX	 ��<�>!t��X��K�|KPLUGG���ǐ��PRCU�B����������Ox��^�SEGF\K:�L�W����Ϟ�����������Q�LAP {ߎ�P#:L^p� ������ >WTOTAL����WUSENU{� i�m>"�RGDISPMMCZ�eR!Cb��@@���OyЛ��ń_�STRING 1�T
�M�MS
�_I�TEM1�  n /!/3/E/W/i/{/ �/�/�/�/�/�/�/?�?/?A?S?e?I�/O SIGNA�L�Tryout Mode��Inp�0Sim�ulated��Out�<OV�ERRx� = 1�00�In c�ycl�5�Prog Abor�3���4Statu�s�	Heart�beat�MH� Faul5G>CAlerHIx?fOxO�O��O�O�O�O�O�O_ ���/_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo8�o�o_WORZ�� �aI_�o�o!3E Wi{����������/�A�S�PO�)Ay��kb��� ����ҏ�����,� >�P�b�t���������pΟ���t�DEV|� ���
�D�V�h�z��� ����¯ԯ���
���.�@�R�d�v�����PALT5]���o�� �����1�C�U�g� yϋϝϯ���������p	��-߯�GRI�� �e�ٿ?ߍߟ߱��� ��������/�A�S� e�w�������S�KR5]	�}���1�C� U�g�y����������� ����	-?Qc<u��PREGž�  !�����/ ASew��������//{=�$�ARG_�`D ?�	���\!��  	�${6	[p(]�p'�{7�)O SBN_CONFIG*@�\+�1�2�!CI�I_SAVE  �{4�!�"O TC�ELLSETUP� 
\*%  O�ME_IO{={<%?MOV_H0%?�+?REP�v?I&U�TOBACK�!�\)�"FRA:\� }?�� �'`@��8�� �;�  �25/11/19� 14:15:52��(�3OEOrOiO�<���O�O�O�O�O__���OA_S_ e_w_�_�_&_�_�_�_ �_oo+o�_Ooaoso �o�o�o4o�o�o�op'9��  �1�_�3_\ATBC�KCTL.TMP DATE.Dļ�������3IN�Iİ�5�%�3MESSAG� �q�!|d �{ODE_D0�&�%�!�O�)��3oPAUSy�!�\+� ,,		�� \%����}��� ��Ïŏ׏���5���1�k�U���y���ş���\�f�TSK  �l��?��0UPD�T ��wd6�6�XWZD_ENB�t�*?�STA�u\!6��N!XIS� UNT� 2\%�!� � 	����v!��ۯƯ ���#��G�2�W�}�n��MET�2���� Ph���d�忈��SCRDCFG �1\%�1 	��%�"ڿ>�P�b� tφϘϿ?�
Q�)+� ������0�Bߩ�f� �ϊߜ߮�������K���G'�1GR��*�J��#�[pNA?0[+	��4 �_ED�p1���� 
 �%{-apEDT-�S:������$60-(�3��
�"�O06���@�  ��-�2 6�R;���O���_��� �#���G�/�3r� O����+������/�4�>b����b��Q�/�5 �
�.���./u�/�/�6f/��/ ����/�/A/S/�/w//�72?�/?�/��[?@�???�?C?/�8�?��KO��'O�O�?�?�OO/�9�O:O_^O����O^_�O�OM_�O/�CR5�m?�_�_ �=�_(oo_�_o�_#�~p�NO_DEL/��!�GE_UNUS�E-��IGALL�OW 1S� �  (*SY�STEM*ɳ	�$SERV_GRpg�ɶ�`f�REG�e�$sɼ�`NUMxz5s#}PMU�`>ɵLAY��ɼ�PMPAL|�pduCYC10on�~lpp~�sULS�Ub$}�rf��cL���tBOXORI�uCUR_�p#}�PMCNV^v��p10�~J�T4D�LIJ���i	*P�ROGRA�dPG_MIp~�����ALz�������B�׏�n$FLUI_RESU�w�
P�@l@o]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y����� h#��LAL_OUT ��k�B�WD_�ABOR�p�o�I�TR_RTN  �+T�:��NONgSTOg�2� �h�CCG_CONFIG S귰T����U�ϟ�e�E_R�IA_I�`2����>�e�FCFGG S�{�+]���_PA�GP 1]����	��B�T�f�%�Cp  ��ނ�Ќ�Ж�Р��Ъ�д�о��Ȫ��҉�܉����މ��  D��D��Ԩ��ݯ��ͽ����� D���	���"	��`D1Z	�9��@�+V?)��e�HE]`l��6�G�_P*�1� ze�ϋ�������������HKPAU�S�1���  �r�G��5�s�Y��� �������������9]oU���O�����+W�CO�LLECT_���������EN�z�2����NDE����c;b�1234567890H6R�a��FXN+S
 Hƿ+S)� ��\����[�� A///0/�/T/f/x/ �/�/�/�/?�/�/? a?,?>?P?�?t?�?�? �?�?�?�?9OO"�a2� ���"IO 1�1X�1ƻO�O�O�O�GTR�	�2mM(8P�I
O�No� �M)ZG�^�I_MORgB!�� ��-�U 	  �Y�_�_�_�_o k�RT�hA"�],G�?0�0��ga�@Kod�A
3�R��#��o�a�bC4  A��qx��� x�@A��z � B�эB�эCo  @�b��@��A:d�
�aI�*$�m�aT_D�EFŁ %�%�7_Rb�&pINUS���F���gtKEY_�TBL  �����` �	
��� !"#$%�&'()*+,-�./Q:;<=>�?@ABC)pGH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������,���͓���������������������������������耇����������������������]A�pLCKpp|\ɋpppSTA��et_AUTO_D�OQ��f�INDx	َ�R_T1��T23�`�M��h�XC� 22v�r��8
SONY �XC-56�o�a}�|`�@���
b} $PА���HR5'SԟR�57���Aff�A]�o� K����� ��ʯܯ�� ���6� H�#�l�~�Y�����B\�TRL(pLETE�0�#�T_SCR�EEN �_kcscc�UM��MMENU 1&~�  <�� @Xϡe7�aϖχs� ���ϩϻ������>� �'�M߆�]�o߼ߓ� ���������:��#� p�G�Y��}����� ����$����Z�1�C� i���y��������� ����V-?�c u����
�� @)vM_�� �����*/// 9/r/I/[/�//�/�/ �/�/�/&?�/?\?RL��_MANUALo�*�DBPQWR�F���DBG_ERRL�.p'&ˮA �e?�?ON�1NU�MLIMT��@d��epDBPXWO_RK 1(&��?�sO�O�O�O�O@]DBwTB_ձ )�=Աc!Q�dy1DB__AWAY�3�a�GCP �b=��EBR_AL1@ُRB�2Yn�ⵕ`�8_�0� 1*�U�AU`
bO�_�d�_�_�H�_M�ISր[@|�`�SONTIM߷���d�f[Y
�upSMOTNEN�DtoTRECOR�D 10&� �<�_�SG�O��a�o �[R�o�o�o�o�h ,�oP�ot��/ E�=�a�(�:� L��p�������ʏ ܏�]����6���Z� l�~�������#�؟G� ��� �2���V�şa� 韞���¯ԯC���g� 񯋯@�R�d�v�寚� ����п?����χ� <�'Ͻ�r�ῖϨϺ� Q�����_�߃�8�J� \���	ߒ�߶�%��� ������4��X����|����!�RTO�LERENCTB��eR*PL�͜0C�SS_CNSTC�Y 21SI�`��cR��+�=�O�e� s��������������� '=K]o���DEVICE 22� �F�� ��
.@Rd�v�_��HNDGDg 3��@Cz�_LS 24�� �//*/</N/`/����PARAM �5|YLR�5r$��SLAVE 6���_CFG 7��/r#dMC:�\��L%04d.'CSVq/5@c?�26R�A >3CHF0�A�_r.Q?�?�'�r&�v2�1�?�9�1X@�JP��3�>cQ�A��,RC_OUT �8��Av/_SG�N 9re[b���mE20-N�OV-25 07�:50A0va1}9ZE14:16A0�� [sr��I�Ar.�@RA@��S�Þ�j���A�N�#VERSI�ON EJ�V4.0.1�\E�FLOGIC 1�:� 	�8�w`)Y�19]RPROG_ENBPh�YSWULSg �R_ACCLIMf���#��SWRSTJN�P2eZcvaQMOb\�1�"�TINIT ;��reva �VOPTι  ?	f�R
 	R575r#VC`74Hi6Ih7Ig#50mh�Dsb2Id�8��oW&dTO  �2m�O�oVV�PDE�X�WdMB� sP�ATH AEJA�\�oQc��HC�P_CLNTID� ?�F�# ��;n���IAG_�GRP 2@�)� xa 	 �E�  F?h� Fx E?`�rD���{�p���Ĺ|����A�/�Cf�J0yJ0Y�dC�J0q�B�i���ymp4m5� 7890123�456���W�p� � A�ffA��=qA�>0хA��HA�>0��ƀ��Ac������1@�>4�p>0���A���,��A0B4�|� �t�2h�1
���(�A��A�
=A��B���A��
A�Q�A��������j�����j!�i0��{+A�Z�̶��Z�>0}����A�ր������h�z��������6�EG�A@�>0:�RA5Z�/�)ր#F�Z� b��P����*�<�6��Pz�AJƀY�?�9p�A3\)�A,��A&�� �����������ȯ6�}cF�]��AW��UP��J��C<Z�u4��-Z�%G�� �0�B�T�6���� ��>�P�ڿ$�rϘ�v� ����X�jϴ��(�� L�^���n�b�pĂQ��ݑi������=�
�==�G���>��Ĝ���7����8��b��7�7y����@ʏ\��p�$�M@�A�h>0/�A��<i���<xn;=�R�=s��=x�<�=�~Z�;7��|�<'��>� �?+ƨC�  <(�U�2w 4����懙����y\�� ? �������6�H�h ��T�~���������������?)7L?S;�F$�/�Y���4G���
�PA1��i�L*�x�A��X�j�|��q����������%��ED  E� ? Eh� DQX�:���1< �0�p����3q�m/�4/:"�yK- #/|/�/y/�/�/�/�/��/�|CT_CON�FIG /v��S�Deg��5�qSTBF_TTS�W
qYP3�@�St�1c6@MAU�P�f_BMSW_CF�$0B�{  	�/JO�CVIEWw0C�=����	OO-O ?OQOcO�R�?�O�O�O �O�O�OuO
__._@_ R_d_�O�_�_�_�_�_ �_�_�_o*o<oNo`o roo�o�o�o�o�o�o o&8J\n� ��������"�4�F�X�j�|��<R%C�3D@Մ2!��� ���؏���1� �U��i4SBL_FAULT E���8o�GPMSKY7��0�TDIAG F�(9�1�	UD�1: 6789012345ߒ58�P�/�-�?�Q�c�u� ��������ϯ���0�)�;�� M��
���

���6TRECP��ʚ
ؔʿ� ����"�4�F�X�j� |ώϠϲ��������π��0�W�i�fߍ�U�MP_OPTIO1NY0{���TR�2Z3:���PMEX5���Y_TEMP  È�3B�}0����A����UNI�0[5�Ѥ6YN_B�RK G�?�2E�DIT_��ENT� 1H��  �,&FGF _�1v�2�&PRO�Gm�� &P�ICKUP���&E���52���(�� L�3�[���i������� ���� ��$6Z A~ew���� ��2VhOЌs��L0EMGDI_STA��,1��A�NC�1I�; �4�&//w�
w�d^߀/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?��O#O5OGOUI m!UO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_]J 
Oo&o8oJodOno�o �o�o�o�o�o�o�o "4FXj|�� ����o��0� B�\of�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�T�J�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ��� � 2��^�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� �����*�<�V�`� r����������� ��&�8�J�\�n��� �������������� "4N�Xj|�� �����0 BTfx���� ����//,/F8/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?��? O O$O>/P/ZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_�?�?�_
oo.oHO Rodovo�o�o�o�o�o �o�o*<N` r����4o�_� ��&�@oJ�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ������8� B�T�f�x��������� ү�����,�>�P� b�t���������֟Ŀ ���0�&�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ�ο�������� :�D�V�h�z���� ��������
��.�@� R�d�v����������� ����2�<N` r������� &8J\n� ��������/ *4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?� �?�?�?O"/O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�?�_�_�_ o O,O6oHoZolo~o�o �o�o�o�o�o�o  2DVhz���_ �_���
�$o.�@� R�d�v���������Џ ����*�<�N�`� r�������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘ߲������� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� �߼����������  2DVhz��� ����
.@ Rdv������� ��/*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?��?�?�?�?/O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�?�_�_ �_�_�?�_o,o>oPo boto�o�o�o�o�o�o �o(:L^p ��_�����_o �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z����� ԟ� �
��.�@� R�d�v���������Я �����*�<�N�`� r�쟞�����̿޿�� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߖ��� �����������0� B�T�f�x������ ��������,�>�P� b�t���|��������� ��(:L^p ������� �$6HZl�� ��$ENETMO�DE 1J���  ����������R�ROR_PROG %�%��/)��TABLE  ���T/f/x/�'��SEV_NUM� �  ���� �_AUT�O_ENB  ����_NO�! �K���" W *� 0� 0� 0	� 0� +� ?+?=?�$HIS�#���+_ALM 1L�� ��� <��+>?�?�?�?�?OOrB?_�"�   ���!�YJ�TCP_VER !��! /$O$EXTL�OG_REQZ69��)�CSIZ�O�D�STK�I�%�~�BTOL  ��{Dzb2�A �D_BWD9@P�&:Q��#SDI(Q M��>S���?[STEPP_b_�|P�OP_DO�O�F�DR_GRP 19N��!d 	TO�_���P�������glpw��qŗ�?�I ���%f�S 7oHm2okoVo�ozo�o �o�o�o�o�o1z�A�c#A���>�ք>��>~8~
 E���� Uq8�SC�"�����xC`}dC�{�N�B�{���}@UUT1�UT��Z��ss��wsM�O�HcEP]��O��#M�˵�/KA��I�?wpя�o�:6:N=���9-��I���,' k�� �o'������B�-�_+�FEATURE �O��:P��Handlin?gTool p����Englis�h Dictio�naryv�4D ;Ste�ardp�x��Analog I�/O����gle �Shiftßut�o Softwa�re Updat�e�matic ?Backupt���ground E�diti�v�Cam�era��FCn?rRndIm�R��ommon ca?lib UIM�u��n4���Monit�or��trn�Re�liabאu�DH�CPi�Īata ?Acquis��ũ?iagnos����߫ocument? Viewe��ǧ�ual Chec�k Safety���y�hancedh��u�^�s1�FrE��w�xt. DIO� ��fi���en]db�Err��L������s��r���� �)Ps�FCTN M�enuJ�vã��T�P In�fac��x�G-�p Ma�sk Exc^�g���HT!�Prox�y Sv2�P�ig�h-Speb�Sk�ih�Q����mmuwnic�ons�ȃur��گ��$�c�onnect 2��ncr#�str�u��t�KAREL Cmd. LK��uaM� �Run-;Ti��Env��밯el +�s�S�/Wv�Licen�seD�1���Boo�k(System�)s�MACROs�,~�/Offse�ސ��H����د��M�R�����Mech/Stop\�t����"��i��ڛ��xb�������odؐwit#ch#����.��I�Optm[���]�f�il1���g�ǅ�ulti-TC�7�t�PCM fun�����o��E�����Re�giz�r����ri�*�F��)���Num� Sel��D��� Adju��?�l�ښ}�tatu%��,��x�RDM Rob�ot��scoveL����em�М�n��|����Servo���6�u�SNPX b�B�ߞSN!�Clix)�8ےLibr��DXe� ��j $o_�=t�ssag��y��m@ ��r�m@/I|"ͱMILIB�~�P Firm��:�P�Acc.�6��TPTXԯ�el�n����m����o�rquؐimul�a��K�uu=�Pa�;��-���W�&\�e3v.��riB�M�USB por[t ��iP��a*��%nexcept�b�����%��h�VC"��r����V��f"�w%jq+SK SC�G�/SUIr�Web Pl���.�� 4d�\�(�߶&�/;7�Grid��pla�y5=� �O7R]".�����-2000i�C/165M���l�arm Caus�e/��ed��As�cii\�k�Loa9d1��:Upl�0P�ycא&�0��O����RA����)y�NR�TLHz�Onh�e Helh���#����#� �z1tr��64MB DRAM]O��CFRO�OB�ell��s�sh�A	_W�cz�U��p�-\t%yאsV�Lt'�s�.s�maiC�NU������qiEL�@Sup"��%��P��A�cro����j}4	<U��Quest�g3miC9q&rtA���r��l�ju�o�o�o�o �o�o�o -$6P Z�~����� ��)� �2�L�V��� z����������� %��.�H�R��v��� ����������!�� *�D�N�{�r������� ���ޯ���&�@� J�w�n���������� ڿ���"�<�F�s� j�|ϩϠϲ������� ���8�B�o�f�x� �ߜ߮��������� �4�>�k�b�t��� �����������0� :�g�^�p��������� ����	 ,6c Zl������ �(2_Vh ������/� 
/$/./[/R/d/�/�/ �/�/�/�/�/�/? ? *?W?N?`?�?�?�?�? �?�?�?�?OO&OSO JO\O�O�O�O�O�O�O �O�O�O_"_O_F_X_ �_|_�_�_�_�_�_�_ �_ooKoBoTo�oxo �o�o�o�o�o�o�o G>P}t�� �������C� :�L�y�p��������� �܏���?�6�H� u�l�~��������؟ ���;�2�D�q�h� z�������ݯԯ� � 
�7�.�@�m�d�v��� ����ٿп����3� *�<�i�`�rϟϖϨ� ���������/�&�8� e�\�nߛߒߤ����� ������+�"�4�a�X� j������������ ��'��0�]�T�f��� ��������������# ,YPb��� �����( UL^����� ���//$/Q/H/ Z/�/~/�/�/�/�/�/ �/?? ?M?D?V?�? z?�?�?�?�?�?�?O 
OOIO@OROOvO�O �O�O�O�O�O___ E_<_N_{_r_�_�_�_ �_�_�_oooAo8o Jowono�o�o�o�o�o �o�o=4Fs j|������ ��9�0�B�o�f�x� ������ȏҏ����� 5�,�>�k�b�t����� ��ğΟ����1�(� :�g�^�p��������� ʯ��� �-�$�6�c� Z�l���������ƿ� ���)� �2�_�V�h� �όϞϸ��������� %��.�[�R�dߑ߈� �ߴ߾�������!�� *�W�N�`����� ����������&�S� J�\������������� ����"OFX �|�������KB  H552?vf21lR78k{50lJ614l�ATUP�545z�6lVCAMlwCRI�UIF��28�NREx5�2�R63wSC�HlDOCV &C�SUx869�0^�EIOC�4k�R69�ESET��J7�MAS�KlPRXY�7.lOCO�(3�kX� ��53C&H�(�LCH�&OPLGz�0�&MHCR�&]S&7MCS�0�'{55�MDSWp7v�'OP�'MPR�&p �&L �PCM��R0�7� �00�75�1�51�80�P�RS'69�&FR�D�RMCNl9=3�SNBA'�'/SHLBHFMjG �c82�HTC�T�MILxC&TPA�[&TPTX�FEL�;F00C'8��wJ�95�TUT�'9�5�&UEC�&UF]R�VCC7XO?6wVIP�FCSC�F�5 IlWEB�H�TT�R6'CG��WIGrWIPGS��VRC�FH7v6�6�R7r'R�:2��&R�*4�&�P�R�64wNVD&Du0&gFIhCLI�8��CMS[&x`�S�TY[WTO�NNn�&ORS?6OL�hWENDxLBWS�hwSLM&FVR[% G*<N`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R� d�v���������Џ�����*�<�N� � H552�P�j�21p�R78�o�50p�J614�p�ATUP��54�5��6p�VCAM�p�CRI�UIFv��28�NRE���52ߚR63�S{CHp�DOCV`�wCSU��869���0��EIOC0�4�o�R69ߚESE�T��ޛJ7ޛMA{SKp�PRXY�]7p�OCO�3���o�젟���53��H�m�LCH�OPL�G��0O�MHCR��S��MCS��0��55��MDSW� �>�OP>�MPR�?�L�/�����PCM�R0~�젯�̰o�[51ϛ51��0Ϛ�PRS߫69/�F{RD�RMCNp�{93��SNBA@�^n�SHLB@�Mn�tL��2��HTC���TMIL����TP�A��TPTX��EL/�̰��8�����wJ95�TUT?��95/�UEC�U�FR�VCC�O�ߺVIP��CSCt��}�Ip�WEB���HTT��R6>�C�G��IG��IPGmS�RC��H7~�[66ϚR7ΫR��2O�R}�4/�\�wR64�NVDߪ�D0��F��CLI_�ΛCMS��, ���STY��TO��N�N/�ORSߺOL�>END��L��S�}SLMߪFVR ��O���
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� ������������0� B�T�f�x������ ��������,�>�P� b�t������������� ��(:L^p �������  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o �o�o�o�o�o0 BTfx���� �����,�>�P� b�t���������Ώ��@���(�:�L�X��STDR�LANGt�o����� ����ϟ����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�e�w߉߸�߭߿�RBTs�OPTN���� ��$�6�DPNr�N�`�r���������� K�� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~�������� 2D9�9N�$FEAT�_ADD ?	����{�  	K��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n�nDEMO O{?   K�� �߽������� ��)� V�M�_�y����� ��������%�R�I� [�u������������ ��!NEWq {������ JASmw� �����/// F/=/O/i/s/�/�/�/ �/�/�/???B?9? K?e?o?�?�?�?�?�? �?O�?O>O5OGOaO kO�O�O�O�O�O�O_ �O_:_1_C_]_g_�_ �_�_�_�_�_ o�_	o 6o-o?oYoco�o�o�o �o�o�o�o�o2) ;U_����� ����.�%�7�Q� [����������Ǐ� ���*�!�3�M�W��� {�������ß���� &��/�I�S���w��� ����������"�� +�E�O�|�s������� ���߿���'�A� K�x�oρϮϥϷ��� ������#�=�G�t� k�}ߪߡ߳������� ���9�C�p�g�y� �����������	� �5�?�l�c�u����� ��������1 ;h_q���� ��
-7d [m������ /�/)/3/`/W/i/ �/�/�/�/�/�/?�/ ?%?/?\?S?e?�?�? �?�?�?�?�?�?O!O +OXOOOaO�O�O�O�O �O�O�O�O__'_T_ K_]_�_�_�_�_�_�_ �_�_�_o#oPoGoYo �o}o�o�o�o�o�o�o �oLCU�y �������� �H�?�Q�~�u����� ���������D� ;�M�z�q��������� �ݟ�	��@�7�I� v�m���������ٯ ���<�3�E�r�i� {�������޿տ�� �8�/�A�n�e�wϤ� �ϭ����������4� +�=�j�a�sߠߗߩ� ���������0�'�9� f�]�o�������� ������,�#�5�b�Y� k��������������� ��(1^Ug� �������$ -ZQc��� ����� //)/ V/M/_/�/�/�/�/�/ �/�/�/??%?R?I? [?�??�?�?�?�?�? �?OO!ONOEOWO�O {O�O�O�O�O�O�O_ __J_A_S_�_w_�_ �_�_�_�_�_ooo Fo=oOo|oso�o�o�o �o�o�oB9 Kxo����� ����>�5�G�t� k�}�������͏׏� ���:�1�C�p�g�y� ������ɟӟ ���	� 6�-�?�l�c�u����� ��ůϯ����2�)� ;�h�_�q��������� ˿����.�%�7�d� [�mϚϑϣϽ����� ����*�!�3�`�W�i� �ߍߟ߹��������� &��/�\�S�e��� ����������"�� +�X�O�a��������� ��������'T K]������ ��#PGY �}������ ///L/C/U/�/y/ �/�/�/�/�/�/?	? ?H???Q?~?u?�?�? �?�?�?�?OOODO ;OMOzOqO�O�O�O�O �O�O
___@_7_I_�v_m_�]   �X�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q����� ����%�7�I�[� m��������Ǐُ� ���!�3�E�W�i�{� ������ß՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߡ߳��������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� �Ͽ���������+��=�O�a�s߅ߗ�  �ؒѳ����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W�Pi�{ߍߝ����� �����������#�5� G�Y�k�}������ ��������1�C�U� g�y������������� ��	-?Qcu ������� );M_q�� �����//%/ 7/I/[/m//�/�/�/ �/�/�/�/?!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�o�o#5 GYk}���� �����1�C�U� g�y���������ӏ� ��	��-�?�Q�c�u� ��������ϟ��� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_�W_i_{_�_�Y�$F�EAT_DEMO�IN  �T���P��P�TIND�EX�[�Qy�PI�LECOMP �P���a��R�U�PSETU�P2 Qe~b�  N :a��S_AP2BCK� 1Ri  #�)�Xno}k%do�o�P`�o�o�Uco�o �o�o)R�ov ��;�_��� *��N�`������� 7���ޏm����&�8� Ǐ\�돀���!���E� ڟ�{����4�ßA� j��������įS�� w�����B�ѯf�x� ���+���O�Ϳ���� ϩ�>�P�߿t�Ϙ� ��9���]���ߓ�(� ��L���Y߂�ߦ�5� ����k� ��$�6��� Z���~����C��� g������2���V�h� ��������Q���u� 
��@��d��q�iH`PLo 2>a`*.VR��Y *�V>�(� PCFoY OFR6:Z�*�NT�P�����,�P�E/'*.F�v/X	�d/�,q2/�/V+STM�/ �/���/'=�/K?V+H?~?7l?)?;?�?W*GIF�?O5��?�?�?TOW*JPG ^O�O5tO1OCO�OO#JS�O_Y �C�O��O%
JavaS�cript7_bOC�S(_�_6|_9_ %�Cascadi�ng Style Sheets�_�- 
ARGNAMOE.DT�_M0�\�_�_Q.d?o�_>.`DISP*5oo�0�o�oQe�a�ooo
�TPEINS.X3ML�o�o:\�o�&aCustom ToolbarG�viPASSWOR�D�oKFRS:�\�I %Pa�ssword Config�&� ��J��n������ 3�ȏW������"��� F�Տ�|����/��� ֟e������0���T� �x������=�үa� s����,���%�b�� �������K��o�� ϥ�:�ɿ^������ #ϸ�Gϱ���}�ߡ� 6�H���l��ϐߢ�1� ��U���yߋ� ��D� ��=�z�	��-����� c�����.���R��� v�����;���_��� ��*��N`��� ��I�m� �8�\�U�! �E��{/�4/ F/�j/��////�/ S/�/w/�/?�/B?�/ f?x??�?+?�?�?a? �?�?O�?�?PO�?tO OmO�O9O�O]O�O_ �O(_�OL_^_�O�__ �_5_G_�_k_ o�_�_ 6o�_Zo�_~o�oo�o Co�o�oyo�o2�o �oh�o���Q �u
���@��d� v����)���M�_�� ������N�ݏr�� ����7�̟[������&���J�ٟ럀�c���$FILE_DG�BCK 1R���m���� < �)
S�UMMARY.DyG��6�MD:�����B�Diag� Summary����
CONSLOG��ׯ�B�����Console� log���	T�PACCNx�ݿ%�ſ��TP A�ccountin����FR6:I�PKDMP.ZI	P6�:�
Nχ����Exceptio�n��<��MEMCHECK��_������Memory� Data�c��9YF)	FTP�u�f���j����m�ment TBD���c�L =�)�ETHERNET���4�������E�thernet ~��figura����}�DCSVRF���m�ߘ��%�]� verify� all��e�M{+�X�DIFF��pv��� �%��diff�����]�CHG01����`����5�����*f`�2�����&1������g�3� �<�`VTR�NDIAG.LS����.!�� ~�nostic/�e�T6a)UPDATES.t�Z7�FRS:\�r��Upda�tes List��4�PSRBWLOD.CM�6�������PS_RO�BOWEL��
�>HADOW$	��/�Shad�ow Changses�/F�*qx"NOTIb�/�/:?��Notifi�c?��/d�+@AG ��?<��?`��?�?� O�?3OEO�?iO�?�O �O.O�ORO�O�O�O_ �OA_�ON_w__�_*_ �_�_`_�_�_o+o�_ Oo�_so�oo�o8o�o \o�o�o'�oK] �o���F�j ���5��Y��f� �����B�׏�x�� ��1�C�ҏg������� ,���P��t����� ?�Οc�u����(��� ϯ^�󯂯�)���M� ܯq� �~���6�˿Z� �ϐ�%ϴ�I�[�� �ϣϵ�D���h��� ��
�3���W���{ߍ� ߱�@�����v��� /�A���e��߉��� ��N���r�����=� ��a�s����&����� \�������"K�� o����4�X� ��#�GY�} �0��f�� /1/�U/�y/�// �/>/�/�/t/	?�/-? �/:?c?�/�??�?�? L?�?p?OO�?;O�? _OqO O�O$O�OHO�O �O~O_�O7_I_�Om_ �O�_�_2_�_V_�_�_ �_!o�_Eo�_Ro{o
o �o.o�o�odo�o�o /�oS�ow�� <�`���+�� O�a���������J� ߏn�����9�ȏ]���j���u��$FI�LE_FRSPRT  ��}�������MDONLY 1�R��u� 
 ��)MD:_V�DAEXTP.Z�ZZ��K�"�1��6%NO Ba�ck file <��u�S�6(��� ���p���ݯ"���� %�7�Ư[����� � ��D�ٿ�z�Ϟ�3� ¿@�i�����ϱ��� R���v��߬�A��� e�w�ߛ�*߿�N��� �߄���=�O���s� ���8���\����~��VISBCKژ|đ�*.VD�|N���FR:\��ION\DATA�\9�����Vision VDO� z������������� ��-R��v�� ;�_���*� N`��7� �m/�&/8/�\/ ��//!/�/E/�/�/ �/?�/4?�/E?j?�/ �??�?�?S?�?w?O�?�?BO��LUI_�CONFIG �S��0�MK '$ +Cߖ{���O��O�O�O�O�OY�@|x4O6_H_Z_l_~_�\ $_�_�_�_�_�_�_
o /oAoSoeowoo�o�o �o�o�o�o�o+= Oas
���� ����'�9�K�]� o��������ɏۏ� ���#�5�G�Y�k�� ������şן韀�� �1�C�U��f����� ����ӯj���	��-� ?�Q��u��������� Ͽf����)�;�M� �qσϕϧϹ���b� ����%�7�I���m� ߑߣߵ���^����� �!�3�E���i�{�� ���H��������� /���S�e�w������� D�������+�� Oas���@� ��'�K] o���<��� �/#/�G/Y/k/}/ �/�/8/�/�/�/�/? �/?C?U?g?y?�?"? �?�?�?�?�?	O�?-O ?OQOcOuO�OO�O�O �O�O�O_�O)_;_M_ __q_�__�_�_�_�_ �_o�_%o7oIo[omo oo�o�o�o�o�o�o��hp|�$FL�UI_DATA �T���.q��a tRESULT 2U.u�Wp �T��/wizard�/guided/�steps/Expert	��� ������0�B��P��Conti�nue with{ GkpanceP� ��������ӏ���	���-�?�Q� r-�q.up�0 �`�`p�0s/q���bpsS�۟����#� 5�G�Y�k�}�����`� �oȯگ����"�4� F�X�j�|���������肟������rip ypğ*�<�N�`�rτ� �ϨϺ������ϯ�� &�8�J�\�n߀ߒߤ� ���������߽�Ͽ��󿱑��tpTimeUS/DST� ���������������0�B�Y�Disably�w������� ��������+=*Or�`8�*�0<�N�`�r�24y�� �&8J\n ��Q�c����� /"/4/F/X/j/|/�/ �/_q����asq?Region�/2? D?V?h?z?�?�?�?�?��?�?U�America� O2ODOVO hOzO�O�O�O�O�O�OU��ayl��/0_�/?>rsditor�O�_ �_�_�_�_�_�_oo�(o:oU� Touc�h Panel �oS (recommenmp)Ho�o�o �o�o�o�o�o/A \�_"_�F_X_>jRaccesO� ���!�3�E�W�i��{�����Conn�ect to N?etwork��ӏ ���	��-�?�Q�c�u�����X��/v؟��!�lPInt?roduct?1� C�U�g�y��������� ӯ� �	��-�?�Q� c�u���������Ͽ�� �Ɵ�꟬ �f�xϊϜϮ����� ������,�>���b� t߆ߘߪ߼������� ��(�:�(�0�>����~d�� Pϵ����������!� 3�E�W�i�{���L߱� ��������/A Sew�H�Z�l�~� ���+=Oa s�������� //'/9/K/]/o/�/ �/�/�/�/�/�/�� �2?�Y?k?}?�?�? �?�?�?�?�?OO1O �UOgOyO�O�O�O�O �O�O�O	__-_?_�/ ?"?�_F?�_�_�_�_ �_oo)o;oMo_oqo �oBO�o�o�o�o�o %7I[m� P_�t_��_��!� 3�E�W�i�{������� ÏՏ����/�A� S�e�w���������џ 㟢��(��O�a� s���������ͯ߯� ��'�9���]�o��� ������ɿۿ���� #�5���V��z�<�>� ������������1� C�U�g�yߋ�J����� ������	��-�?�Q� c�u��FϨ�j����� ����)�;�M�_�q� �������������� %7I[m� ��������� 0��Wi{��� ����////�� S/e/w/�/�/�/�/�/ �/�/??+?�4 X?�?D�?�?�?�?�? OO'O9OKO]OoO�O @/�O�O�O�O�O�O_ #_5_G_Y_k_}_<?N? `?r?�_�?�_oo1o CoUogoyo�o�o�o�o �o�O�o	-?Q cu������ �_�_�_&��_M�_�q� ��������ˏݏ�� �%��oI�[�m���� ����ǟٟ����!� 3����x�:����� ïկ�����/�A� S�e�w�6�������ѿ �����+�=�O�a� sυ�D���h��ό��� ��'�9�K�]�o߁� �ߥ߷���������� #�5�G�Y�k�}��� ������������� C�U�g�y��������� ������	-��Q cu������ �)��J�n 0�2�����/ /%/7/I/[/m//> �/�/�/�/�/�/?!? 3?E?W?i?{?:�?^ �?�?�/�?OO/OAO SOeOwO�O�O�O�O�O �/�O__+_=_O_a_ s_�_�_�_�_�_�?�? �?�_$o�?Ko]ooo�o �o�o�o�o�o�o�o #�OGYk}�� ��������_ (ooL�v�8o������ ӏ���	��-�?�Q� c�u�4������ϟ� ���)�;�M�_�q� 0�B�T�f�ȯ���� �%�7�I�[�m���� ����ǿ������!� 3�E�W�i�{ύϟϱ� ���ϔ������ܯA� S�e�w߉ߛ߭߿��� ������ؿ=�O�a� s����������� ��'�����
�l�.� �������������� #5GYk*�|� �����1 CUgy8��\�� ����	//-/?/Q/ c/u/�/�/�/�/�/� �/??)?;?M?_?q? �?�?�?�?�?��?� O�7OIO[OmOO�O �O�O�O�O�O�O_!_ �/E_W_i_{_�_�_�_ �_�_�_�_oo�?>o  Obo$O&o�o�o�o�o �o�o+=Oa s2_������ ��'�9�K�]�o�.o ��Ro��Ə����� #�5�G�Y�k�}����� ��ş������1� C�U�g�y��������� ��ʏ����ڏ?�Q� c�u���������Ͽ� ���֟;�M�_�q� �ϕϧϹ�������� �ү���@�j�,��� �ߵ����������!� 3�E�W�i�(ύ��� ����������/�A� S�e�$�6�H�Z߼�~� ����+=Oa s����z��� '9K]o� ����������/ ��5/G/Y/k/}/�/�/ �/�/�/�/�/?�1? C?U?g?y?�?�?�?�? �?�?�?	OO��� `O"/�O�O�O�O�O�O �O__)_;_M___? p_�_�_�_�_�_�_o o%o7oIo[omo,O�o PO�otO�o�o�o! 3EWi{��� ��o����/�A� S�e�w���������~o ���o��o+�=�O�a� s���������͟ߟ� ���9�K�]�o��� ������ɯۯ���� Џ2��V������� ��ſ׿�����1� C�U�g�&��ϝϯ��� ������	��-�?�Q� c�"���F��ߺ�~��� ����)�;�M�_�q� �����x������ �%�7�I�[�m���� ����t߾ߘ����� 3EWi{��� ������/A Sew����� ��/����4/^/  �/�/�/�/�/�/�/ ??'?9?K?]?�? �?�?�?�?�?�?�?O #O5OGOYO/*/</N/ �Or/�O�O�O__1_ C_U_g_y_�_�_�_n? �_�_�_	oo-o?oQo couo�o�o�o�o|O�O �O�O);M_q �������� �_%�7�I�[�m���� ����Ǐُ�����o �o�oT�{������� ß՟�����/�A� S��d���������ѯ �����+�=�O�a�  ���D���h�Ϳ߿� ��'�9�K�]�oρ� �ϥϷ�ȿ������� #�5�G�Y�k�}ߏߡ� ��r��ߖ��ߺ��1� C�U�g�y������ ������	���-�?�Q� c�u������������� ����&��J� ������� %7I[�� ������/!/ 3/E/W/x/:�/�/ r�/�/�/??/?A? S?e?w?�?�?�?l�? �?�?OO+O=OOOaO sO�O�O�Oh/�/�/�O  _�/'_9_K_]_o_�_ �_�_�_�_�_�_�_�? #o5oGoYoko}o�o�o �o�o�o�o�o�O_�O (R_y���� ���	��-�?�Q� ou���������Ϗ� ���)�;�M� 0B��f˟ݟ�� �%�7�I�[�m���� ��b�ǯٯ����!� 3�E�W�i�{������� p����������/�A� S�e�wωϛϭϿ��� ���ϴ��+�=�O�a� s߅ߗߩ߻������� �¿Կ�H�
�o�� ������������� #�5�G��X�}����� ����������1 CU�v8�\�� ���	-?Q cu������ �//)/;/M/_/q/ �/�/�/f�/��/� ?%?7?I?[?m??�? �?�?�?�?�?�?�!O 3OEOWOiO{O�O�O�O �O�O�O�O�/_�/>_  ?_w_�_�_�_�_�_ �_�_oo+o=oOoO so�o�o�o�o�o�o�o '9K
_l._ ��fo����� #�5�G�Y�k�}����� `oŏ׏�����1� C�U�g�y�����\� �ʟ����-�?�Q� c�u���������ϯ� 󯲏�)�;�M�_�q� ��������˿ݿ￮� ��ҟ�F��m�ϑ� �ϵ����������!� 3�E��i�{ߍߟ߱� ����������/�A�  ��$�6Ϙ�ZϿ��� ������+�=�O�a� s�����V߻������� '9K]o� ��d�v����� #5GYk}�� ������//1/ C/U/g/y/�/�/�/�/ �/�/�/���<?� c?u?�?�?�?�?�?�? �?OO)O;O�LOqO �O�O�O�O�O�O�O_ _%_7_I_?j_,?�_ P?�_�_�_�_�_o!o 3oEoWoio{o�o�o�_ �o�o�o�o/A Sew��Z_�~_ ��_��+�=�O�a� s���������͏ߏ� �o�'�9�K�]�o��� ������ɟ۟ퟬ� �2����k�}����� ��ůׯ�����1� C��g�y��������� ӿ���	��-�?��� `�"��ϖ�Z������� ����)�;�M�_�q� �ߕ�T���������� �%�7�I�[�m��� PϚ�tϾ�����!� 3�E�W�i�{������� ��������/A Sew����� �������:��a s������� //'/9/��]/o/�/ �/�/�/�/�/�/�/? #?5?�*�?N �?�?�?�?�?OO1O COUOgOyO�OJ/�O�O �O�O�O	__-_?_Q_ c_u_�_�_X?j?|?�_ �?oo)o;oMo_oqo �o�o�o�o�o�o�O %7I[m� ������_�_�_ 0��_W�i�{������� ÏՏ�����/��o @�e�w���������џ �����+�=��^�  ���D�����ͯ߯� ��'�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗ�N� ��r��ϖ�����1� C�U�g�yߋߝ߯��� ���ߤ�	��-�?�Q� c�u��������� �����&�����_�q� �������������� %7��[m� ������! 3��T�x�N� ����////A/ S/e/w/�/H�/�/�/ �/�/??+?=?O?a? s?�?D�h�?�?� OO'O9OKO]OoO�O �O�O�O�O�O�/�O_ #_5_G_Y_k_}_�_�_ �_�_�_�?�?�?o.o �?Uogoyo�o�o�o�o �o�o�o	-�OQ cu������ ���)��_�_oo ��Bo����ˏݏ�� �%�7�I�[�m��> ����ǟٟ����!� 3�E�W�i�{���L�^� p�ү������/�A� S�e�w���������ѿ ������+�=�O�a� sυϗϩϻ����Ϟ� ��¯$��K�]�o߁� �ߥ߷���������� #��4�Y�k�}��� ������������1� ��R��v�8ߝ����� ������	-?Q cu������� �);M_q �B��f�����/ /%/7/I/[/m//�/ �/�/�/�/��/?!? 3?E?W?i?{?�?�?�? �?�?��?�O��? SOeOwO�O�O�O�O�O �O�O__+_�/O_a_ s_�_�_�_�_�_�_�_ oo'o�?Ho
Olo~o B_�o�o�o�o�o�o #5GYk}<_� �������1� C�U�g�y�8o�o\o�� Џ�o��	��-�?�Q� c�u���������ϟ� ���)�;�M�_�q� ��������˯��ԏ�� ��"��I�[�m���� ����ǿٿ����!� ��E�W�i�{ύϟϱ� ����������ܯ�  ��t�6��߭߿��� ������+�=�O�a� s�2ϗ��������� ��'�9�K�]�o��� @�R�d��������� #5GYk}�� ������1 CUgy���� �������/��?/Q/ c/u/�/�/�/�/�/�/ �/??�(?M?_?q? �?�?�?�?�?�?�?O O%O�FO/jO,/�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�O�_�_ �_�_�_�_oo/oAo Soeowo6O�oZO�o~O �o�o+=Oa s������_� ��'�9�K�]�o��� ������ɏ�oꏬo� �oҏG�Y�k�}����� ��şן������ C�U�g�y��������� ӯ���	��ڏ<��� `�r�6�������Ͽ� ���)�;�M�_�q� 0��ϧϹ�������� �%�7�I�[�m�,�v� P����߆������!� 3�E�W�i�{���� ���������/�A� S�e�w���������~� �ߢ�����=Oa s������� ��9K]o� �������/ ������h/*�/�/ �/�/�/�/�/??1? C?U?g?&�?�?�?�? �?�?�?	OO-O?OQO cOuO4/F/X/�O|/�O �O__)_;_M___q_ �_�_�_�_x?�_�_o o%o7oIo[omoo�o �o�o�o�O�O�O�O 3EWi{��� ������_�A� S�e�w���������я ������o:��o^�  ��������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�*���N� ��r�׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫�|��� ���Ŀ��;�M�_�q� ������������ ���7�I�[�m���� �������������� 0��Tf*���� ����/A Se$������ ��//+/=/O/a/  jD�/�/z�/�/ ??'?9?K?]?o?�? �?�?�?v�?�?�?O #O5OGOYOkO}O�O�O �Or/�/�/�O
_�/1_ C_U_g_y_�_�_�_�_ �_�_�_	o�?-o?oQo couo�o�o�o�o�o�o �o�O�O�O�O\_ �������� �%�7�I�[�o��� ����Ǐُ����!� 3�E�W�i�(:L�� p՟�����/�A� S�e�w�������l�ѯ �����+�=�O�a� s���������z�����  �'�9�K�]�oρ� �ϥϷ��������Ͼ� �5�G�Y�k�}ߏߡ� �����������̿.� �R��y������ ������	��-�?�Q� c�t������������ ��);M_� �B�f���� %7I[m� ��t����/!/ 3/E/W/i/{/�/�/�/ p�/��/��//?A? S?e?w?�?�?�?�?�? �?�?O�+O=OOOaO sO�O�O�O�O�O�O�O _�/$_�/H_Z_O�_ �_�_�_�_�_�_�_o #o5oGoYoO}o�o�o �o�o�o�o�o1 CU_^_8_��n_ ���	��-�?�Q� c�u�������joϏ� ���)�;�M�_�q� ������f��ԟ�� �%�7�I�[�m���� ����ǯٯ�����!� 3�E�W�i�{������� ÿտ�����ʟܟ� P��wωϛϭϿ��� ������+�=�O�� s߅ߗߩ߻������� ��'�9�K�]��.� @Ϣ�d���������� #�5�G�Y�k�}����� `���������1 CUgy���n� ������-?Q cu������ ���/)/;/M/_/q/ �/�/�/�/�/�/�/? �"?�F?m??�? �?�?�?�?�?�?O!O 3OEOWOh?{O�O�O�O �O�O�O�O__/_A_ S_?t_6?�_Z?�_�_ �_�_oo+o=oOoao so�o�o�ohO�o�o�o '9K]o� ��d_��_��_� #�5�G�Y�k�}����� ��ŏ׏����o�1� C�U�g�y��������� ӟ������<�N� �u���������ϯ� ���)�;�M��q� ��������˿ݿ�� �%�7�I��R�,�v� ��b����������!� 3�E�W�i�{ߍߟ�^� ����������/�A� S�e�w���ZϤ�~� ������+�=�O�a� s��������������� ��'9K]o� ��������������DN�$FM�R2_GRP 1�VL� ��C4  B]� 	  ����E�� �����OHcEP]���O��#M{���KA����?�/��:�6:N�.!9-��6%�A�  �R/d+BH�C`}�dC��N�!B�{�%���/�-އ@UUT�/UT���/?�>���>c��>rа�=ȫ�>i��=���.����:��:���:/:6)�:��~�/s??p?��?�?�?�?�?`_�CFG WmT �?=OOOaOK�NO m
�F0�A �@LRM�_CHKTYP  ] uw-_�ROM�@_MIN\�@���@�� ]X`SSBCXL ��_S1_C_	ETP�_DEF_OW � uXWIR�COM�@i_�$G�ENOVRD_D�O�F�]THR��F d�Ud�T_E�NB�_ �PRA�VCfY�GP ��I_4o�?Xo�qfowo�* ��Q�OUi_m�A��mR�<�@ -�o�o�o6+C�����L_$�Zr%tfq|s���iJ_�PSMTf`�
iyP[t�$HO7STCB1amP�� 	1�&1�1�a�	e}�����ҏ�� ���'�9�K�n�o���	anonymousr�����ğ֟� 0�B�T�1�h���� y���������ӯ��� 	��>�t���c�u��� �������(�*�� ^�;�M�_�qσ�ʯ�� ���������H�Z�7� I�[�m��ƿؿ��� ����2��!�3�E�� V�{��������� ����/�A��ߚ߬� ������������� `�=Oas��� �������\� n���.������ ����/#/5/G/ jk/��/�/�/�/�/ 0BT1?h/�g? y?�?�?�?��?�?�? 	OO>?t/�/cOuO�O �O�O�/??(?*O_ ^?;_M___q_�_�?�_ �_�_�_ _�_HO%o7o�Io[omo��ENT� 1b�k P!\o�o  �p�o �o�o�o2�oV b=��s��� ���@���v�9� ��]�����⏥���� ۏ<���`�#���G�}� ����ޟ���ş&�� 2��[���C���g�ȯ ��쯯��ӯ�F�	��j�-���Q�QUICC0��w���꿭�A1�ǿٿ:ϭ�2;���)ϊ�!ROU�TER��g�y���!?PCJOG�϶��!192.168.0.10��~��CAMPRT+��!�1$�R�9փRT��V�h��ߏdN�AME !�j!�ROBOD���S_CFG 1a�i� �A�uto-star�ted�DFTP�Ob��O�_��*_�� ��������_�/�A� S�v�d�
��������� ���N;�M�_�<s��� S�������� &I�\n� ����O�O�O�O5 "/iF/X/j/|/�/U �/�/�/�/�//�/0? B?T?f?x?�?��� �?	?�?=/O,O>OPO ?tO�O�O�O�O�?aO �O__(_:_L_�?�? �?�?�O�_�?�_�_ o o$o�OHoZolo~o�o �_5o�o�o�o�o  g_y_�_h�o��_� ����o��.�@� R�uv�	�������Џ �);M_a�3�� r�����������ޟ� ��&�I�˟\�n��� ���������!�ϯ5� "�i�F�X�j�|���U� ��Ŀֿ��ϟ�0��B�T�f�x����_ERR c�ڈϘ��PDUSIZ  ��^7����>~��WRD ?)�����  guest����,�>�P�b���SCD�_GROUP 3�d)� -�#�� ��LOA��n��RES��TM�޷ $��T_��E�NB��TTP_A�UTH 1e��� <!iPen�dann�y����.!KAREL�:*y���KC������VISION SET��)� �-!@�.�X��� |�j����������������H�CTRL Kf��b�
��FFF9E3���FRS:D�EFAULT��FANUC W�eb Server�
uH����0��/AS��WR�_CONFIG �g��������IDL_CP�U_PC� �B����� BH�M�IN����GNR_IO������ȭ�NPT_SIM_�DO�+STA�L_SCRN� ��]!TPMOD�NTOL='+�RTY(�
&�L�E��='�ӪOLNK 1h�����/�/��/??'?9?�"MA�STE��)
%O�SLAVE i���h5RAMCAC�HEW?O"ON�O_�CFG�?�#�3UOx(�?�2CYCL�?��5� _ASG 19j���
 ;?>O PObOtO�O�O�O�O�O��O�O__(_C;BN�UM����
�2I�P�?�7RTRY_�CN� ��ʭ29!_�UPD���!��� �2�0�2kw>���_��ЭSDT_IS�OLC  w;����J23_DS�$U-`OBPRsOC�/	%JOG�Ի1lw;<�d9<���?�3[�o"3_?ï���lQ�o &8�o\n���o%hr`��1�_+b�P�0EVo&KANJI_Q0K�
���?MON m��b�yWp���������H�Υ��Sn�lڅ�L$��_L�NRq_��EYLOGGI�N�0�М�a����$LANGUA�GE ��"�� ����LG�Ro�I�! ��xJ�భp�������'0Ȥ�;�|�j ;��
�(UT1:\ȏ� �!�3�E�\��i�{�������ï�(�_����LN_DISP pw?ߘ�o��o&�OC["�Dz���A��OGBO_OK q��d�0e�桳�Xޜ׿ �����cJy��5�S�e	��������Ϩ����_BU�FF 1r�-��2��ϲ�m�ϐ �,�Y�P�bߏ߆ߘ� �߼���������(��U�L�^��=���DC�S tKNp=���P̏�Jx9������)���IO 1u�K �_b�� b�r������������� ��&:J\n ���������=�E�TM	nd �k}����� ��//1/C/U/g/ y/�/�/�/�/�/u�@�SEV�P6�<TYP	nZ;?M?_?�-�qRS�P/��éR�FL 1vK��P����?�?�?	OO-O�?Op?TPC�	o*2>o�NGNAM6d~��v���UPS.�GI�U���U�A_LO{ADS`G %6��%PICKUP�1LO8\MAXUALRMNW$\XP�A'_PR�T�P ��Q�PC1�w��9��x]XPt`P 2x^[W ���	*1͐��P�|_Nt�R�_ �_�_(o��oWoBo{o ^opo�o�o�o�o�o �o/S6H�t �������+� � �a�L���p����� ��ߏʏ����9�$� ]�H�����v�����۟ ��П���5� �Y�k� N���z��������ԯ ���1�C�&�g�R��� n��������п	�����?�*�c�WDBG?DEF ylE���jQl�~�_LDXD�ISA�@kK;�ME�MO_AP�@E {?lK
 �� J������"�4�F�X��j�PISC 1z
lImP�UϷ��T�π��P����*�ύ�_MSTR {�-~M�SCD 1|���"���������� ����>�)�b�M��� q������������� (L7p[m� ������" H3lW�{�� ���/�2//V/ A/z/e/�/�/�/�/�/ �/�/??@?+?=?v? a?�?�?�?�?�?�?�? OO<O'O`OKO�OoO��O>�MKCFG �}\�v_�SLTAWRM_�B~�W�B��P�B��$_,TUPM�ETPU��;c���d�ND�PADCO�LFU��Q^CMNT�g_ ZUU� �\�^SQ�_�TZUP�OSCF�W�^PgRPM�_�YSTeP{1�\� 4@�@<#�
Ua�AUeeo sgQosouo�o�o�o�o �o�o�o5)kM�_�����qZQS�ING_CHK � j_$MODA�QS����K�N�D�EV 	\�	�MC:E�HSIZ�E�͜@��TAS�K %\�%$1�23456789� ��ą�TRIGw 1�\� l\�%m���C��9��SF��YP�$�'���EM_INF 1��	W��`)�AT&FV0E0�F���)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ�����H�=�̑1�e���Am���P�����ݯ� ���ǟٟ ���n�!���ɯ��ȿ {�쿧��"�	�F��� �|�/�A�S���Ͽ�� ��1�����T��x� _ߜ߮�a��߅ϗϩ� ��,���P��a��9� ��e������������ :���������G�� ����������6 Zl��C�U�g�y� ��� WD��h�#y���>�NIwTOR�PG ?Y��   	EX�EC1�C"2(3�(4(5(Հ&7*(8(9�C"� p$
"p$"p$""p$." p$:"p$F"p$R"p$^"�p$j"p#2w(2�(2��(2�(2�(2�(2��(2�(2�(2�(3�w(3�(3"�R_�GRP_SV 1݄�� (�q�H�V�>�c=u�q������?Y<@�@����_Da���3ION�_DB�@���A/  �@Q4�E-MK��@4���N 0�E
4�-ud1k��O�O�O�A�PL_NAME �!�U�@�!�Default �Personal�ity (fro�m FD)PB>PR�R2�1 1�L?68L@P�A�P
 d�R_-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_oqo�o�oTC2_�o�o �o�o,>PbTB<�o����� ��
��.�@�R��H�ED  ��\  �  ��  ��0A� W B��T���eB���� g �����0B���p���  CT@C�T@P Ez � E�� E�` E�τ;߈΅ҁ��τZ�䏖π�  E�� �΁΁[�@����ЃTӀA#��׀�2�:�� F�2�N�ޅ�2��~�
��g��7��΁� �:�����2�2�ʝޕޘɂ3��.��΀Dځ�D���*� �1��~����~�0�@���F�:���/3�Jт�3�(����c��:�ڀ�E	˘Em���1�ޥ��ޥ
��� U�g�y��� ������ӿ���	��-�F�,�R�d�v����w�E��QEw:U\��  ���0  ������TBd��w��������$�����J6��RG'4� � W%�I߂ߔ�  hتߠ�A��A��������ߧ�����º����B�0��K�[�TB�	`��ߎ���q�:��oAPI������RG ������B�C��IP�|�0 ��P(� @�?�0j�N�?xT@j�TA@�6I��jH��;�	lz�	�  ���pX�0�H@���X �� � �, ����0K�l,K����K��2KI�+�KG0�K �Uq�E��-3��0@6@ t��@�X@I��V��{��N�����
��}?v����S ���j %��
=�ô�ڀ�h�!�b��澺����a�fҶ��T@�1 V�HA!�2H��Z~�xz�	'�� � �I�� �  ����t�:�È�ß�=����@���T�/}T��!/iOAd/�  'z&G{ ?���V� R�UC� B��C0C� �Bڀ�!�JT@���Cp����� `02C�B ��6P@5��:5TAD΀y�_?u߃?n?�?l�?�05f@�`�2��	 ٠T�"�5 �� ��:Ɓ���{�?�ff05�O*O�? k�_O�qK8���O�J?Y��Ҁv�:(���EP��H�9����,#?3�33O$�E�;�x�5;��0;�i�;�du;�t�<!�	CO���z�T�z��?ff�f?�?&tPB�@��A#�Q@�o[�U#)�"oQ ���7j��_h��_XW�� IOo	oBo-ofoQo�o�uo�o�o�o�o%(��F'0�o �oD�_e��Y7�3xEC� �_.���� �9� $�]�H���l�����B/ ؏����Z �~G��� k�}�����@_��ȟb� ����
�C�.���'0cA�l��}� C>�`��:�5U���� �8�� ���ĩ��W$�C�d��` #Ca!��뤿���V ܢ.��bC�@_;C9�B�A�Q�>�V�È�����Y�uü��
q�C���Q���hQ�A��B=�
?h����#���W���ÈK�B/�
=�������=&�K�=�J�6XK�r#H��Y
H}��A��1&�L�j�LK����H:��HK��b�t�	bL ��2J��8H���H+UZBu&����������!� �E�0�i�T�yߟߊ� �߮��������/�� ,�e�P��t����� �������+��O�:� s�^������������� �� 9$IoZ �~������ �5 YD}h��������G�y�// C�a{�>// Ĉ��Q/X/OCVF�y/�/�=�<�/����K�/�/� 
E�/�/�/??zҰ(ұ�_�hA?��A��r5��N���b?t?��3lC�8�?�?�2�ⷺ?�?��t�.3��}��?�<k���q'�3�JJMIRO@@OvOdO�O�LåP2R	P�N���OH?_0+__O_:[�U_\_��_�_�\{�_�_�1  fU�_�_oo=o (oao_ڏ�o�o�o�k�Ͼo�o�o�o{)�Z   ( 5�o�<6�r�����x  2 wE%p��E[@�w�N���Bw�k�w�C%�`�t���@E/@� ��;�]�o�������Ĩ�������9�(ԁԇ9���mQ9�rYa��ɫ
 $� ��������ϟ��� �)�;�M�_�q�Ⱥ������;I�v��$MSKCFMA�P  E� �va�]�֮���ONREL  ��E���@��E�XCFENB�
8����FNC���JOGOVLIM��d���d��KE�Y�_�h�_P�AN�z�v���RU�NO�{�SFSP�DTY�@����S�IGN��T1M�OTQ����_C�E_GRP 1�E��\RoV�Jo zό��tvϷ�n��ϒ� �����5���*�k�"� �ߡ�X���|����߲� ����U��y��r� ��f�������	�����QZ_EDIT�����TCOM_C_FG 1���l��d�v���
D�_AR�C_��E>�T_?MN_MOD	0����UAP_C�PL��"�NOCH�ECK ?�� �E+�!3E Wi{��������/ܫNO_WAIT_L�l9�$�NTL����zc��_ERR.�s2����A� �����+���"/4/� ��O���| G �J��/�1<��|0?Z��/�/\�q.��PARAM�����&o/!?cW��L? =�p345?678901f?x? �:a?�?�?�?�?�?O`�?'O9OKbW�kO�}L?�O�ODRD�SP����OFFSET_CAR/����FDIS�O�CS;_A��ARK�:��OPEN_FIL�EP��:���OPTION_IOp����[PM_PRG ;%��%$*�_�^�7SWO#P�4��#� �U���RFΠ �Q��P�G�Q	 �+��Q��Q����@RG_DS�BL  �����d�`o�ARIENTkTO��Q�C�[������@UT_SIM_DcW�����@�V�@LCT � �6��T���iQ�g��a�_PEX��_�dR[AT�� d��d>�@UP ��nr�9��WiO��y��$�"2-ÈL�68L@P�c
 d�O��� �*�<�N�`�r����� ����̏ޏ����&�8�J��(2�z����� ��ԟ���
���# i�F�X�j�|�������@į֯�����(O4�a��D�� � ��  �� A��  BI�/�B���s9�H=���  ��E�� BJI�pI�Ȅ`�a#`�P Ez  E��� E�` EE���;������ቴ�Z�������  �E���������@V������T��Aݸ���ر����� �챀ɘ����ر8�ر�!Ģ�Ա����ر�� @Ŭ����쵄͘ŘȂ������ر��D����D��ر������ ��8�H���8���ż���� ���X�/�ǋ���(U�t������f��E	��`�EmYԀ���Ƙ��ͼ����Ř� �!�3�E�W�i�{����������F�����0�:��/�	9H�m���c�D ����������P�P��M�'4 � �W%<�/ �0:dZ
At�A�m����wa�*��t���B`���80�P$:	`�NHZl�:��o�a����i@Г��t�pO=p1��+[�+v���t60�+dP( �@�ծ!�!!?�(C���u�  ;��	l�"	 ` ����pX�M0.�q �X� � � �,� ��"80H��9�H�H���H`�H^yH�R+!h]��/4�,80C�`B�I����C44A ?5�9|]�t��
=Ç`��D1(?:?L?9Bz��Βa#am�$?9p��?�#`9!�3.��=�-��/A�F86O4	'� � TB�I� �  ���.
=���8xO�K�2@�O�@ �>,a�O;K,b�4�?��?'@N�P"_  'fP:T1a0B@�2�`�2u?G_Y_ 3�  ϥ�C*�&���վ.`�P21B� �V�P�U��A�U#aD��3o/Ao�,oeoPo�05�p��`�bUA	 S٠�R�e �  � �:��R"�Q�4�?��ff���o�ozo !%/{8+�E�Sz?Y��4!Xj(+��uP�x�i�!�#�$^�C?333Q$��1�;�x5;��0�;�i;�du�;�t�<!���/�6$�C8"��?fff?�@?&�2�]d@��A{#H�@�o[P� '��R-�J&Zg(%��&' ���l$܏Ǐ �� $��H�3�l�~�i��� ����؟ß��s�����X��V��E���� 쟝������������ ��?�*�c�N� _�� \�R/�޿<��x�)� ;�M�_��tφ� Ϲπ��������ύ �PA1�*��;� C��a�p���u����?�M�����߼�^'�gD��W��C�" �` !C�2)�ж�Կ�Ш��L�@I�`^���bC@_;C9��BA�Q��>V��È�����Y�u�ü��
/������Q��hQ�A��B=�
?�h�è�� ���W��ÈK��B/
=�����Ɗ=��K�=��J6XK�r�#H�Y
H}���A�1��L��jLK����H:��HK� �2�	bL� �2J��8H���H+UZBu�߅������ ��������'7 ]H�l���� ���#G2k V�z����� /�1//U/@/R/�/ v/�/�/�/�/�/�/? -??Q?<?u?`?�?�? �?�?�?�?�?OO;O &O_OJOoO�O�O�O�I�Gϭ�O�O C��a9��O Ĉ��<__CVF�7_>_����_�@��K<�_�_� 
E�_�_�x_�_x�(xѳ_ʙh�_�q��0e�E��N�� o2o��3l�C�Lo^olb���xo�o�t�.3��}�o�lk���q'�3�JJ�m �i�o4"XF|��%P�rP�~������o�����{� ��S�>�c�{c�r��a  fU��N�׏ �������R�@�v�d��|��������̛)Z̟ޟ  ( 5�-�����B��0�f�T�����  2� E%p��E[-@��N���B5�)і5�C��2Ј�@ _���"�4�F�X�i����������ɿۿP�㾡����x�+�����|ԇ�
  �E�W�i�{ύϟϱ� ����������/߆�����tkI�v��$PARAM_MENU ?�e��  �DEFPU�LS�\	WAI�TTMOUT���RCV�� S�HELL_WRK�.$CUR_ST�YL�P��OP9T���PTB�����C��R_DECSN��{uN�H�Z�l�� ������������%�� �2�D�m�h�SSR�EL_ID  ��e�q�|�USE_PROG %w�q%i���}�CCR�����q���_HOSoT !w�!��#��T�p��?�A{��_TIM�E�Ҏ���h�GD�EBUG��w�}�G�INP_FLMS��P��TR��P+GA  ����CH��TYPE
t���h�b��� ���	///(/Q/ L/^/p/�/�/�/�/�/ �/�/ ?)?$?6?H?q? l?~?�?�?�?�?�?O��?O OIO�WOR�D ?	w�
 �	PR� �MsAIE��SU�ƄCTEb �EH	�ԑBCOL��I�O�FTRACECToL 1��e��W �p�p_|S�FDT Q��e�JPPD � zsW_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��S_���� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������� �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ����������1�C��M��$PGTRA�CELEN  �N�  ���M��c�_UP ��������~�  ��c�_�CFG ����|�M������r�������  �����DEFSP/D ���L�u���c�IN��TROL �����8���:�PE_CONF�I������������c�LI�D�㞲�	��GR�P 1�u�� lN�C% � ��l�M�A��;H�N������A�  D	�� ��r�	\M�d`��	!	�������������; ´tV?Bw �~h�z����"�Bz�/A+� <}�<�oFB|��� �^�!/�1/W/B/"��z|#�/M�
l/�/ \/�/�/�/?�/+?? O?:?s?^?p?�?�?�?�?�?��)M�)
�V7.10bet�a1�� @��@�A&�ff��*AC  kC� �<CDk���S@C�LD�@ DĠ Dr� ��cBH� 
���C5<B� N�?�  �ACCpO�E������MXM�O|CAp���`�O
__._�����KNOW_M � ����SV {�������/�_�_�_�?�_�_��_o����M��sZt��:B	��<A��� o�o�\id+ `�`2��@
�+A�
��e�o�l����MR*��QmT�
�xCM�Cf�#�8J{��S�T��1 1����P4���x$u��� �������%� �)�n�M�_������� ڏ��ˏ���F�%�7�I�hw2s|]a�M�G�<������3������Пhw4����#�hw5@�R�d�v�hwA6������ɯhw7���
��hw89�K�]��o�hwMADo� ��厕OVLD  ����o"�htPARNUM  v{��#�isSCH޹ ��
u�>���|��UPD>��Q�ό�_CMP_G`o����L�'����ER_CHK���ib֌��RSpU_��_#MO�g�y�_cߋ��_RES_Grp���
�B��������� �"�S�F�w�j��� �������ɼ�ә��������� �?�D� ��?�_�~����Ӓ��� ������������� 8�;@�Ӌ�[z<��V 1�vu�Ѿ]a@b��y�T?HR_INR�Х��/b��d�MASS6� ZMN�-�MON_QUEUE �vu^V���AU��N��U@�N=f}END��ߜ�EXE����BE���}OPTIO���ۀPROGR�AM %`%��d�~TASK�_I��OCFG� �`R�T/� D�ATAJc��+@�&2�f�/	??-? ??�/c?u?�?�?�?V?��?�?�?O�.INFOJc��-�o�?]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_@�_�_�_�_ G,D��,c ��!��K_�!���)LNfG�!2��k X,	}	J�=���\o���i$3�Xa�i�i��g_EDIT ���/�o�_� WE�RFL��esRG�ADJ ��jA�  #u?��/u�v�a�vuO�?��j�!<xa��LF%����h�oEsf�Q2�Qw>B	Hw�l���^q>�㻎A��t$��*�/� **�:����#�?�D��X�S����q]�D� �p�}�K���[�m��� �����Ǐُ���� ��3�E�s�i�{����� ��ߟ՟�a���K� A�S�ͯw��������� 9����#��+���O� a�������ϻ�Ϳ�� ��}�'�9�g�]�o� �ϓϥ�������U��� �?�5�G���k�}߫� �߳�-�������� ��C�U��y����� ��������q��-�[� Q�c��������������	�/h�V�z ���}�y�AwPREF ��Qz��
uIOORITY'�f�qMPDSP
!�jyr�oUTr&�svOD�UCTo!�j��vOG�P_TG��`t"�j�TOEN�T 1��k (�!AF_INE��+/6'!tc�p6/^-!ud�M/�.!icmXu/�~�XYJs��l;��a)� +��/�/�`��/%?5? Q?8?u?\?n?�?�?�? �?�?O�?)OOMO_O	*�Js�Qyyr��O��O�s>�%�%B+�/5��O_�t��x��~Asr,  �G�QO_a_s_�_�e��0�8JrqPORT_NUM���`�eq_C?ARTREP�`�n�3`SKSTA� �jLGS( ��k�ss�`Un?othing�_ko�}o�o/`TEMPG ���o&S`�_a_seiban��o�4X C|g����� ���	�B�-�f�Q� v����������Ϗ� �,��)�b�M���q� ����Ο��ޟ��(� �L�7�p�[�������ʯ��iVERS�Ix�� �disabled���SAVE ���	2670H�721���{�!`�O}����/�� 	׸H�(	� �ce� F�X�j�|ϊ�5̲��ϵ,?�_� 1�
�+h���B�������)URGE_�ENB�|��QW�FD�DO��R�W�$ e��Q�ZWRUP�_DELAY ���^X�R_HOT %M��O��v��R_NORMAL������)���SEM�I�.�m�'QSKKIP����W��x߯ ��ۯ���������+� �O�a�s�9������� ��������9K ]#m����� ���5GY }k��������/1/C/���$R�BTIFf�lRC_VTMOUg�%��a DCR��¾�� ���8�+K�k�Ed���A��C����3=C���Q���lqk�?|���D2	����?3;�x5;���0;�i;��du;�t�<!���?��	?r?�= K_�?�?�?�?�?OO�%O7OIO[OmO�WRD�IO_TYPE � ��c?yOEFP�OS1 1�G��Pxֿ�J��`?__ =_ʿa_�O�_ _�_�_ V_�_z_o�_'o9o�_ �_ o�olo�o@o�odo �o�o�o#�oG�ok ��<N��� ��1��U��R��� &���J�ӏn���	��������Q�<�u��OOS/2 1Ħ��O,��f��b�����A3 1Š���ğ��|�g�|���S4 1�5��G�Y������5���S5 1�ʯܯ�(�𦿑�ʿH�S6 1�_�q�����;�&�_�>ݿS7 1������R��ϻ���r�S8 1ʉϛϭ���e��P߉��SMASK 1˖O �@����N��XNO�O���<��AMOTEh �K��,�_CFG ��3�~���BPL_�RANG/�k/m�O�WER ��������SM_DRY�PRG %��%�0����TART �Θ���UME_�PRO����B��_�EXEC_ENB�  X5s)GSP�D�]�e��!t�TD�B����RM����I�A_OPTION�&� u#'�MT_���T��1�w!a O�BOT_ISOL�C��b�_�N�AME ���1��IOB_ORD_NUM ?����AH72�1  X4�@Ȯj �
Z��PC�_TIME�'o)x�a S232L�1���)8LTEA�CH PENDA1N� H��P=/���Mainte�nance CoKns�>`"Z��No Use P>�Q�����{!
NPO�������CH_Lf��x�	y!~D/!UD1:�/zF/R��VAIL������'�SR + ����g�J-�R_INTVAL������*0���)V�_DATA_GR�P 2���*!*�D0P{ߝ?w��?�9 ���?�7�?O O6O$O ZOHOjOlO~O�O�O�O �O�O�O __0_V_D_ z_h_�_�_�_�_�_�_ �_o
o@o.odoRo�o vo�o�o�o�o�o�o *:<N�r� ����� �&�� J�8�n�\��������� ���ڏ���4�"�X��F�h���|���'��$�SAF_DO_PULS� (�C!*�ܑN̐CAN�����L SC���+��(+����W���`�P������ �? d�v���������M�������*�<�(JC#ע2e���de�‱�2n�G� @�f㬿��п⾔��� ��0��_ @#T���?�Q�c�~p�T D��p� �ϫϽ��������� )�;�M�_�q߃ߕߧ���/%�������)#��=;W�o$$p55�%
�t��D�i� ء<��� � �;
<�4�$��� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew���������� �//0/S�\/n/ �/�/�/�/�/�/�/�/1@/��0M��X�� O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o�CoUogoyo�o�o �o�o�o�oP/	- ?Qcu��?25 <?ע����!�3� E�W�i�{��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p�0������������ ��� ��$�6�H�Z� l�~�������ƿؿ�����ۯ%�R�\Ɨ����K�!�	�1234567�8��h!B�!ܺ�tա٠ /0��������
��.� @�R�X�گ{ߍߟ߱� ����������/�A� S�e�w����j��� ������)�;�M�_� q�����������������BH (:L ^p�������� $6H��;�jT~��� ����/ /2/D/�V/h/z/�/�/��D� �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?��O&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_Oj_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o [_�o�o�o�o, >Pbt�������ɤ���'���oL�^�p���C�z  Aз�  W �}�2͢���} }�
ɇ�  	į�����X�+�9�>�����;��㏈�������П �����*�<�N�`� r���������̯ޯm� ��&�8�J�\�n��� ������ȿڿ���π"�4�F�X�jτ��b�;�ׁ��<���$�SCR_GRP �1�+�8+��  � ��a� ��	 ���� ������<�����v���p!��H߀����~E�D�` D�W���Ë�E�f�R-�2000iC/1�65F 5678�90ـ��ـR�C65 ���
O1234�����G  ɋ������X���%���f���E����+�	��|�����������H���]��������@�3�E�����a �@�����ȟ���h�����BǙ�B��  B�33B� ������A��G  @�`6��@{ЎF  ?L�^��H���o!
��F@ F�`������ ���
C.g ��4f�}���B��V/�+// O/:/L/�/p/�/�/�/ �/�/W�:o�1�7D?���ˀA?v?�b^@L�6�X�|?�3Bh6 �?����7�� ��%��O�A{���H1C_�[�<@f�0B��a ROyO�O�JgAp�H�O�O�O P�B(�B�O_"_�/F_1_�j_tV��EL_DE�FAULT  ~/����`��SHOTSTR��]=A�RMIPOWERFL  ��x�U���QWFDO�V� �U�RRVENT 1�������U L!DU�M_EIPt_9h��j!AF_IN�E�PWo�!FT$-o�nMo�o!���o� ��o�o!RPC_MAIN�o��h��oB	sVIS��i�1�!TMP�pPU�@id}��!
PMON_�PROXY�Cfe �&��r�<mf�r��!RDM_SR�Vs�@iga���!�R��ڏAhh��
�!%
pM=�=li��V�!RLSYN���r�}�8E���!gROS,oɜ�4����!
CE�pMT'COM�Cfkݟ:�{!	�CONS;��Bgl)���!�WOASRC��Cfmu�vү!�USBӯAhn����oB���� !�k���W���{�ؿ������WRVICE_�KL ?%k �(%SVCPR#G1�K�5�2K�P�":�3s�x�:�4�Ϡ�":�5����:�6����:�7��:���[�V�	9c�h�7�Տ��:� =ϸ�:�e���:���� :���0�:���X�:�� ��:�-ߨ�:�U���:� }���b��� �b���H� b���p�b���b�F� ��b�n���b���b� ��8b���`b��� ��6���:�!�3�� ��@+dO� s�����/� *//N/9/r/]/�/�/ �/�/�/�/�/?�/8? J?5?n?Y?�?}?�?�? �?�?�?O�?4OOXO CO|OgO�O�O�O�O�O �O�O_	_B_-_T_x_�c_�_�_DEV �i�MC�:���*��TGR�P 2�e� /��bx 	� 
 ,`�_o�o Ho/oloSoeo�o�o�o �o�o�o�o DV =za��o�� �
��.��R�d�K� ��o��������ɏ� �*�<�#�`��U��� M�����ޟ�ן��� 8�J�1�n�U������� ȯ���ӯ�"�y�F� X�?�|�c�������ֿ ������0��T�;� xϊ�qϮϕ�����;� ߿�,�>�%�b�I߆� ��߼ߣ�������� ��:�!�^�p�W���� ����������$�� H�/�l�~�e������� �������� V ��z�s���� �
�.RdK �o�����/ /o</�`/r/Y/�/ }/�/�/�/�/�/?�/ ?J?1?n?U?�?�?�? �?/�?�?�?"O	OFO XO?O|OcO�O�O�O�O �O�O_�O0__T_;_�M_�_�Sd ԑV	 x_�_�_�_�_	o�_-o�<k%�<oao�S���za&aze�o�g�o �o�o�o�o yNo3 vi�o`N�r�� �� �D�8�&� \�J���n�����ݏ ������4�"�X�F� |������l�֟h�� ���0��T���{��� D�����ү������ ,�n�S������t��� ��ο��޿�F�+�j� ��^�Lς�pϦϔ��� ���ߺ��϶�$�Z� H�~�lߢ�����ߒ� ������ �V�D�z� �ߡ���j��������� �
��R���y���B� ������������Z� ��Q��*�r�� ���2V�J �Z�n���
 �.�"//F/4/V/ |/j/�/��//�/�/ �/??B?0?R?x?�/ �?�/h?�?�?�?�?O O>O�?eOwO.OPO*O �O�O�O�O�O_XO=_ |O_p_^_�_�_�_�_ �_�_0_oT_�_Ho6o loZo|o~o�o�oo�o ,o�o D2hV x�o�o���� �
�@�.�d����� T���P�Ώ���� <�~�c���,������� ��ʟ�ޟ�V�;�z� �n�\���������Ư �.��R�ܯF�4�j� X���|�����ٿ뿢� Ŀ���B�0�f�Tϊ� ̿���z��������� �>�,�bߤω���R� �ߪ����������:� |�a��*����� ������B�h�9�x�� l�Z���~�������� ��>���2��BhV �z�����
 �.>dR�� ��x��/�*/ /:/`/��/�P/�/ �/�/�/?�/&?h/M? _??8??�?�?�?�? �?�?@?%Od?�?XOFO hOjO|O�O�O�OO�O <O�O0__T_B_d_f_ x_�_�O�__�_o�_ ,ooPo>o`o�_�_�o �_�o�o�o�o( L�os�o<�8� �� ��$�fK�� �~�l�������؏Ə ��>�#�b��V�D�z� h�������ԟ���:� ğ.��R�@�v�d��� ܟ��ӯ��������*� �N�<�r�����دb� ̿��ܿ޿�&��J� ��qϰ�:Ϥϒ��϶� ������"�d�I߈�� |�jߠߎ��߲���*� P�!�`���T�B�x�f� ��������&��� ��*�P�>�t�b����� ���������& L:p�����`� ��� "H� o�8����� �/P5/G/� /� h/�/�/�/�/�/(/? L/�/@?.?P?R?d?�? �?�? ?�?$?�?OO <O*OLONO`O�O�?�O �?�O�O�O__8_&_ H_�O�O�_�On_�_�_ �_�_o�_4ov_[o�_ $o�o o�o�o�o�o�o No3ro�ofT� x����&�J �>�,�b�P���t��� ����"�����:� (�^�L���ď����r� ��n�ܟ� �6�$�Z� ������J�����įƯ د���2�t�Y���"� ��z�������¿Կ
� L�1�p���d�Rψ�v� �Ϛϼ��8�	�H��� <�*�`�N߄�rߨ��� ��ߘ����8�&� \�J���ߧ���p��� �������4�"�X��� ���H����������� ��
0r�W�� � x�����8 /��P�t� ���4�(// 8/:/L/�/p/�/��/ /�/ ?�/$??4?6? H?~?�/�?�/n?�?�? �?�? OO0O�?�?}O �?VO�O�O�O�O�O�O _^OC_�O_v__�_ �_�_�_�_�_6_oZ_ �_No<oro`o�o�o�o �oo�o2o�o&J 8n\~��o�
 ���"��F�4�j� �����Z�|�V�ď�� ���B���i���2� �������������� \�A���
�t�b����� �������4��X�� L�:�p�^���������  ��0�ʿ$��H�6� l�Zϐ�ҿ�������� |��� ��D�2�hߪ� ����X��߰������� �
�@��g��0�� �����������Z� ?�~��r�`������� ���� ������� 8n\������ �� "4j X����~�� /�//0/f/��/ �V/�/�/�/�/?�/ ?n/�/e?�/>?�?�? �?�?�?�?OF?+Oj? �?^O�?nO�O�O�O�O �OO_BO�O6_$_Z_ H_j_�_~_�_�O�__ �_o�_2o oVoDofo �o�_�o�_|o�o�o
 �o.R�oy�B d>�����*��lQ���q�$SE�RV_MAIL � �u���v�O�UTPUT���v�RV 2���  �� (�"�`��z�TOP1�0 2�Ɖ d �-�?�Q�c�u� ��������ϟ��� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�����YPE����FZN_CFG ����� ���Z�G�RP 2�k�W� ,B   A��~!�D;� B����  B4!��RB21��HELLd���U�ـڏ����#�%RSR#�$�6�o�Zߓ�~� �ߢ����������5�� �Y�D�}����  �q������,���� !���������2!�d�����L���HK 1��� ����� ������������%  2Dmhz��������OMM ����$��FTOV_ENB��΁U�d��OW_REG_U�IDx�IMIOFWDL���y/WAITAE���Ȥ��e̈́�TI�Me���VA����y_UNIT�@&U�LC^TR�YeU�z�MO�N_ALIAS k?eՀheK� �/�/�/�/�*�/�/? ?0?�/T?f?x?�?�? G?�?�?�?�?O�?,O >OPObOtOO�O�O�O �OyO�O__(_:_�O ^_p_�_�_�_Q_�_�_ �_ oo�_6oHoZolo ~o)o�o�o�o�o�o�o  2D�ohz� ��[���
�� �@�R�d�v�!����� ��Џ⏍���*�<� N���r���������e� ޟ���&�џJ�\� n���+�����ȯگ� ���"�4�F�X��|� ������Ŀo����� �ɿ/�T�f�xϊ�5� ���������ϡ��,� >�P�b�߆ߘߪ߼� ��y�����(���L� ^�p���?������ �� ���$�6�H�Z�l� ���������q�����  2��Vhz� �I����
� .@Rdv!�� ��{�//*/</��`/r/�/�/�/S#��$SMON_DE�FPROG &�����!� &*SYS�TEM*�/�'�L�@�$REC�ALL ?}�)� ( �}4co�py frs:o�rderfil.�dat virt�:\tmpbac�k\=>127.�0W01:2372��/s?�?�?  }+�.2mdb:*.*�C?U;Z?�?�?O�8/x.4:\�?8@R>�?PoO�O�O�40.Ea6O HO_A_O�O__�3-? ??�?b_t_�_�_�?F_ �?a_�_oo)O�OMO �_po�o�o�O8oJo�O��o �Utpdisc 0R^�o�o�j|��Ytpc?onn 0 7I [���#_5_�_Y_ j�|����_�_N��_� ���o1o�oUof�x� ���o�o@������ ��-�?�ȏb�t����� ��F�Ϗa����)� ��M�߯p�������8�@J�ݟ� �ϥ�-���:prog_1.;tp��empȯܿ�m�ϑϤ�..�ickup;�O�^���� �&�8���ܯm�ߑ� ����Q�Z������"� 4�ǿX�i�{��� C�ֿ������0�B� T�e�w����߮�I��� ����,��P� s����;��`����
xyzrate 61 �@��n����.�R�72.31.3=2��65968N `�//��.x� ��l/~/�/��q9/@K/]/�/ ??%1[���/�/�/p?�?�?'����18308 @L?^?�?OO&�./ �7�?�?mOO�O�/�+ DOVO�O�O_�.���@�>�Op_�_�_'�1�π?_�;`_�_oo(�7.�@��_8ovo�oo �ŵ�Po�2^o�o�%��$SNPX_�ASG 2�����9q�o  0%�%��a  ?�*vPA�RAM �9u�Cq �	O{P�%�%�dx�t��,pOFT_KB_?CFG  %�?u�)sOPIN_SI�M  9{�r�
��.�8�,pRVN�ORDY_DO � �u�uJ�QS�TP_DSB�~��r��!{SR �>9y � &�zя�"�&vTOP_O�N_ERRW��P_TN 9u+���C�RIN�G_PRM�i�V�CNT_GP 2��9u�qFpx 	 ����%�s�����П%w�VDZ�RP 1��y�p��5����� /�A�S�z�w������� ��ѯ�����@�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥ��������� ���#�5�G�Y�kߒ� �ߡ߳���������� �1�X�U�g�y��� ������������-� ?�Q�c�u��������� ������);M _q������ �%7Ipm ������� /6/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaO�O�O�O�O�O�O��O�PRG_CO7UNT�v�+�Y'ENB@�UM0S�t�=__UPD 1�>��T  
�O�b �_�_�_�_�_�_�_o o)o;odo_oqo�o�o �o�o�o�o�o< 7I[���� �����!�3�\� W�i�{�������Ï� ����4�/�A�S�|� w�����ğ��џ�� ��+�T�O�a�s��� �������߯��,� '�9�K�t�o������� ��ɿۿ����#�L� G�Y�kϔϏϡϳ��π������$��1��L_INFO 1�uY[P ��@Tߘ߃���ߧ���OOA���H��о3����� �3Z�5A��@[j�����y¿��CGE�LYS�DEBUGPvP��H�d^Y&�SP_PwASSUB?8�LOG �uU]Q  H����Q�  �ZQH�UD1:\d�X�e�_MPCj�uU����uQ��� uQ��SAV �m�$Q��؍��G���SV��TEM_TIM�E 1�m��P+ 0HЎHԍ����z�SKMEM  �uU Q��  �H�%��H�� �PH����H���H�"R��[PAT�0P;	��H��
�Hс�����ZQ^�� W*:	U� j|��������//0/B/T/�� Z//�/�/�/�/�/�/ �/?!?3?E?W?i?{?��?�?�?�?�?eQT1?SVGUNSpPU�'^U��0ASK_OPTIONP�uUZQ$Q
A_DI�G�1_&EBC2_G_RP 2�uY���4lOH�@7 C��C�<�BCCFG ��YK\���N` �O��_�O_C_._g_ R_�_v_�_�_�_�_�_ 	o�_-ooQo<ouo`o �o�o�o�o�o�o�o;MH�8|g9 ��'����� *��J�D�R�x�f� ���������ҏ��� �>�,�b�P���t��� ������Ο��(�� L�:�\�^�p�����wp ��̯������2� � B�h�V�������~�Կ ¿����
�,�.�@� v�dϚψϾϬ����� ����<�*�`�N߄� rߔߖߨ�����︯ �,�J�\�n��ߒ�� ������������4� "�X�F�|�j������� ��������B0 Rxf����� ���>,b� z����L�� /(//L/^/p/>/�/ �/�/�/�/�/�/�/ ? 6?$?Z?H?~?l?�?�? �?�?�?�?�? OODO 2OTOVOhO�O�O�Ox �O�O
__._�OR_@_ b_�_v_�_�_�_�_�_ �_oo<o*oLoNo`o �o�o�o�o�o�o�o 8&\J�n� ������"��O :�L�j�|�������� �֏��0���T� B�x�f����������� �����>�,�b�P� r����������ί� ���(�^�L���8� ����ʿܿ�l�� � "�H�6�l�~ϐ�^ϴ� ������������ � V�D�z�hߞߌ��߰� �������
�@�.�d� R�t�v����� ���*�<�N���r�`���������������$�TBCSG_GR�P 2����  ���� 
 ?�   'K5oYk@������������d0
?���	 HD z�@$>����BH��CPD�)��L��n>g���2cCP�Rdvp��Cj�� 'B�#B����YxG!7fff
)C�(/*/ ��S)?�.'��( �%�/�/�/?9???d?�?�;?�P#����	V3.00~�2	rc65�3	*�0�4���?�64wW4pf9 @�=�O  � �� �|?UO\C��J2������\OhHCFG ����J��(O�N��O_Z��_A_,_ e_P_�_t_�_�_�_�_ �_o�_+ooOo:oso ^o�o�o�o�o�o�o�o  9$6oZ� ~���r'���� �+��;�a�L���p� ����͏ߏ����'� �K�6�[��������� ������ʟ ��$�� H�6�l�Z�|�����Ư ���د���� �2� h�V���z�����Կ¿ �
���.��R�d�$� |ώ�8Ϯ��Ͼ����� ��<�*�L�r߄ߖ� Tߦߨߺ������&� 8�J��n�\���� ����������4�"� X�F�h���|������� ������
TB xf������ �� 2�bPr t�����// (/:/�^/L/�/p/�/ �/�/�/�/�/? ?6? $?Z?H?~?l?�?�?�? �?�?�?�? OODO2O TOzOhO�O�O�O�O�O �O�O�O
_@_._d_R_ �_�_D�_�_�_�_o �_*ooNo<o^o`oro �o�o�o�o�o�o& J\n�:�� �����"��F� 4�j�X�z�|���ď�� �֏���0��@�f� T���x�����ҟ��� ���,��_D�V�h�� ������ί����� �:�L�^�p�.����� ����ȿ� ��̿޿ H�6�l�Zϐ�~ϴϢ� ���������2� �V� D�f�h�z߰ߞ����� �����
�,�R�@�v� d������z����� ����<�*�`�N���r� �������������� 8&\J���� p�����4" XF|j���� ���//B/0/R/ T/f/�/�/�/�/�/�/ ?�/?>?,?b?��� �?�?H?v?�?�?O�? (OOLO:OpO�O�O�O dO�O�O�O�O�O$_6_ H_Z__~_l_�_�_�_ �_�_�_�_ ooDo2o hoVo�ozo�o�o�o�o �o
�o.>@R �v������ �?�0�B��r�`��� ����������ޏ�&� 8�J��n�\�������Π�  ܐ�� �������A��*SYSTEM*ܐ�V9.0055 �!�1/31/20�17 A p � �D�TBJ�OP_GRP_T�   $ $�F2MGNT�$�MINF2]�CO_MP_SWT�ܐ�D�PARAMN��� $$MR_MAX_TRQ]��R_STAL��B�RK��VEL��N�OLD��A_LOKAD��D۬��_Z�AJ�AV ��������̢Z�D�D�D:+�D:�PTHJ�����ST���,���N�=�DYN_FRCx �ʤ��R_ACͷ�R_DE�LON�G �J����³T� �SP1,�f�SPU3,�4,�5,�6,ĥ7,�8]�x�JJ�c ��s��EL3��  	��f���A�SYM_}��� �����2��SH�ORTMO_SC`ã���b��SH��; ��UMA�����Z���Z�_CYC_?ID 	#�+�_E3�0�f�0�C�0��PAYܢ
�2J_�UP�NGn�LW�y�w�kه�Z�INE�RTIA_VIB���؞���V_U�NIT����f�R_F2J����������������%����RJ_S��L���c�]��HVAà��$H�Z�z�AXO���$�FLEX������TM�HR_TAB�LE S���E}N�� $DIˠ���DO��u���CFGN� )0U���I��A\������_TI � �ME� u���� � � k�MEN��$�u���T��PT+И� �B�L��NU��$CEN:�H�c�W�T9��[� $DUM�MY1C�$PS�_OVERFLO�Wܐ$����F;LA��YPE�¸��K�$GLB_T�������C���T�ORQCTR�� � X $DgEBU@�K�ST���  $SBR���M21_V��� T$SV_ERb��O-�1CL��>ACTIO����GL��EWN� �4 $M�$Y*]�Z]�W|P�g��A���w�^Ub� U�N� .�$�GIF.�}$b ��\� N�	� Lm �,�}$F�,�E�NEARPwLAN��$F�DI��NCw�J�OG_Rޡ 
�u�$JOINT�����MSET.N�  �E��oCONS��
��ONFN�� �$MOU.�?�� LOCK_FOyL���BGLV=��GL�TEST_sXMàoEMPB�)���$U1S8�c O�2 �B�	�n����CENEa" $�KARE��M��T�PDRAe 8$/V�ECLE��/IU��
�HE�TOkOLO�m$VIx#;REP IS3f��&96K���ACHU���{!ONI���29��� I��  �@$RAIL_B�OXE�� RO�BO�?�HOWWAR���!��!OROLM��5A���6SK�"��M�O_�F60! ��G�#0CHN�;��R�S OCN�;SL�ODH0C�O�UW��E�LECTE-Л�$PIP�NODE�"�"�!���[0� ?CORDED����z1��P6 � o D ��OB�T�G�1�����2p,�A��1ADR�ܢ�C�TCH�� 7 ,U�EN���A�_�iDW����ZVWVA�� � > b��P�REV_RT\��$EDIT�FVS�HWR60P��@I)Sv��D-�3���Df�$HEA�D=�r��@M��CK�Ev��CPSPD.VJMP@L��� oRACE��@�^II�SBCH�ANNEw AT'ICKx#��M��o��?SHN�� @P@\QZ��CI�P�V��&��STYcB�!L�O��K?R�RO�� t 
�@GoE%�$�A�= S�!$��O�2�����9P���VSQU2 ,��LO���TERC�G�l��TSDT� � L�33!BDE$�g��Te!��OH�;�F/�IZ�������PR�0���b��0P9U���e_DOh@�XSSK��AXIt�`43�UR_p0��$T� �P'Fb�RgEQ_e 9BET:rQP�@���PF��2�PA�������#l�#�� ��SRJ�lz`��H�� �u���y���u̧�sک �s��u��u��u,���'�Y��K��+�C��9�CJ�%�7�I�[����SSC��  h DS�P���3SP��'�AT�¢��a�PhR��ADD�RESx#B�@SH�IFz�_2CH��#AI��y��TuU��I�� ;�CUSTO[tx�V
�I��ZB�;���*��
�
�RV�1�aN�� \�0�8��Pɜ�a���CX��b^r�ؚ�67��TXS�CREE�2��aTINAT� Y�·�;q;�{� TNQ4 ��A3�p���qBr���@RRO��� �P�����UEDT ���RA��9SUARSM�P�gUNEXd`�����S_�0�^� �3�N��^�;qC���� [2T�UEw���Ds��`GMTɰL�}�q  OE�B�BL_� Wd�� S ��PвO�ܲ�LEk��� ���RwIGH�BRDF�a�CKGRd��T�EX)p��WIDTH�#�@���O���UIC0EY;��! dm �����R� �aBACK��Q�b��J&�FO��1��LAB�q?(�&�Iv�$UR��!����d�,�Hơ O" 8|� _�Ay���-�Rv ��#�'H����Or��#�PIQ�U��<�R��1LUM<�v[�E#RV�1Z d�P
k�5$$�opGE���4fp�)�@LP��dr	Ea`Q)��Q�����آ ��5��6��7��8��_b;��`
�Ԍ��!�S��#�c�USRb% �<�0,�U����F�O���PRIwqmx� *��TRIP�!�m�UN����&� `���e1�e�8�8p2` '��X�.�aG `T40ځLz���OSK���R>p̢��t!�(k}�� �Tư�U���)�)�;�I��һU��OF�F��* Q�O�� 1( ����-) GU3AP��irp��ׁ��x�SUB�R�M ��SRT"�t+0�R@0�cOR� ,'RAU�p-TB	_G��VC�p�,�# �"�1)c$~�=a�#��CW�DRkIV�fEq_VP��@�D9�MY_UBY8��V �)eء>`q��A�!�P_S@	 �kB�M�$gPDEY�dCEX��䣤!�P_�MU3PX�s%�US7Q���` p�Zb}�萐آ[aGl�PAC3INwQ&`RG�`������F��X�uR!E�o�t!ire��X0- ��TAR�G� P<� ��fR�X0.s�5�qY��	t�aRESW&�_A�kpt�`�ON�a�As�{#�rE")�U�P�!kpI@f+HK�R/�P�*~�0�qx ���#EA�P�'�WOR) {%��"MwRCV��0 ���UO�PM) C=�	28��#2REF��-6 6�!j x�hsR ]�:�c1!:c12;�56�/_CRC�+�8�+#�S&��k��a���"��1 ��Rl�Y�5pj��|`OU�W��V�� ,%ہ2-`��Z���`wP.:�tہcRKpSULg`�/h�CO��0eb@�C���C�A�F ѯFE�Cn@L�E`)�E��GE��x>DT2| +:�pqz݀ :�CACH�SLOW1+TAQfFYP��H��SC_LIMIl�FRoXT�qV�;�$HO) b/PC'OMM��O���W`H1���"DԀVP"$4p�R_�f�TZ��XlpP�XWA�UMPjWFAIpPG�$@P�ADDiuIMRE!Ddb�WGP�[�p�pASYNBUFpVRTD�e�d�Q6+�OLt�D_��euWF�P��ETUT�]PQ� �eECCU�VEM�*UrpWVIRCDa�e�c��>�a_DELA��qX���
AG�iRhGXYZR�:�hW8!vsx�#pT� ���"yr��3����LASF�H;1Q�Gqa�4��]QSf`<VN�t/ LEXEU5��\p�Y:�~#FL�I\�cFI�`����KB�#�"?q(�"6d����4=�E��ORD���Qᜓ(B�U7d�_�T����b�OO�;ҥ SFJ���8  f�x�Ah[UR~"SLۀM��#9��[W�J��k3�'a��:��Ç���LIN���X�VR��;����T_�OVRp�
�ZABC<"��v�2��bZ���=��DB�GLV�SL����  �ZMPCEF>�ؐ���.�LNK92
֒i? ЇдQ� �CMCM�C�SC�ART_,�94P_~7� $JJ�D�D�QP�a�Z��f���;2UX�q�UX!Ez���qU���k���������������Z���@ ��ɔ�p	��Y[�D�� Ab��RR`��~�HE
�H��ć��Z���ư|젍�B � Є881���EAKk�0K_SHI��` �RVpF�2��|�C��E�:��Dр������2Iӳ�UD�T�RACE �V���SPHER,��C ,j@'�=�O�#��$TBJO_� �2 ���X�/���k��	J�Q�X�� �	  ���pXm�� ���� �� �,k� �@q�i�	 �D� ��CaD��k�i��������>���� ��<�!a���?�����>L��B� � B��A�L�D�)�^�CQp�D��S����>����~���fff��?�\<���^�&ًC 4Р8���\�D5m�ΣԚ݊�/��2�333<���^�>���>��&�C������k�Cj��~�kߙ����j�;�9bB��*�?8Q��p�P�Hl���|���Y���3��/�A�;��y6��.�>u.�DP���������3��A�/�<Z;u���������& \�N8Ft��: ����5��TnXf�����k�  ��	V�3.00o�rc�65n�* n����)* F� � F�� F�� F�  G�� GX G'�� G;� GR�� Gj` G��� G�| G�� G�� G�8� G�� G�<� H� H�� H��; Ez � E�@ E��� EK F� F[ F�c F�� F�� F�PE"G �� GpU#?h �GV� GnH �G�� G�� �G�( =k�=�+�8�$�ZP0)-?!1k�$3?�  ��V?d:J�'ESTð��X�q��c�s3H�@T��1�X�S�B0k�d897 ��@9d7d8�k��d8d8	d8
d8�d8�5k�d8d8:d8�6RDI�?b��?�?�?�?�?EtDO|O�K�O�O�O�O�N�2SzO`� >J�_�_ �_�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�oi=yP}_a±78y !_3_E_W_OO'O9O`KO]H�2r`� Xūb����p pn@o@�2� ��s��@J�2�BF_�TT1�u`�ԐI�V�ERmCJq_�I�R� 1�; 8$/k����� ��C  ����ȏڏ��� �"�4�F�X�j�|��� ����ğ֟�1����g�B�T�j�x�����A0Is��Ư��MD���Ɯ�  �2�D�V_qIX�j�D�INT��Ģ�D�T�ؿ� Bpas�Ϣ�_TC8τJ�D�$��tφ��R�Q�Ϻω�_�v�@���v0MI_CH�ANU� �� #�D_BGLVLU����u1&�ETHERA�D ?��y��"0���ϒߤ�n8&�oROUT��!Z�!������SNM�ASKn؎S�255.4��2�D�V���v0OOLOFS�_DI0��X�O�RQCTRL !���s%?��T���� 
��.�@�R�d�v��� �������������(��K:os3PE?_DETAILؙ��PGL_CONF�IG �����/cell/�$CID$/grp1s��1�s���\n��� �E���/"/4/ �X/j/|/�/�/�/A/ S/�/�/??0?B?�/ f?x?�?�?�?�?O?�? �?OO,O>O�?�?tO@�O�O�O�O�OB~}cO __(_:_L_^_�q`�_e]�bO�_�_�_�_ oo\O9oKo]ooo�o �o"o�o�o�o�o�o #�oGYk}�� 0������� C�U�g�y�������>� ӏ���	��-���Q� c�u�������:�ϟ� ���)�;�ʟ_�q� ��������H�ݯ�� �%�7�Ư[�m����𣿵�ǿ� �U�ser View� �	}}1234?567890��
� �.�@�R�Z�����z���޹2�W����π������uχ��3 ��d�v߈ߚ߬߾���ߍ�4S��*�<�N� `�r��ߓ��5��� ������&���G���6�������������9�����7o�4FX@j|������8# ��0B�c�i lCamera���@����/�BE� ,/>/P.��j/|/�/�/�/�/��  ��ɗ ?&?8?J?\?n?/�? �?�??�?�?�?O"O4O[��R��?�O�O �O�O�O�O�?�O_"_ mOF_X_j_|_�_�_GO YG�7_�_�_o"o4o Fo�Ojo|o�o�_�o�o �o�o�o�_YG�+�o Zl~���[o� ��G �2�D�V�h� z�!�n��ď֏� �����B�T�f��� ��������ҟ䟋�YG "	{�0�B�T�f�x��� 1�����ү����� ,�>�P���YG�	篜� ����ҿ������,� >ω�b�tφϘϪϼ�c�u�9H����!�3� E�W���hߍߟ�Fϰ߀��������/�
	�0��j�|���� ��k��������0�B� T�f�x���1�C�� .�����+=�� as������� �����+�Oa s���P��� </'/9/K/]/o/ P�cK/�/�/�/�/? ?�9?K?]?�/�?�? �?�?�?�?�/�%�[r? 'O9OKO]OoO�O(?�O �O�OO�O�O_#_5_ G_�?�%;{�O�_�_�_ �_�_�_�Oo#o5o�_ Yoko}o�o�o�oZ_�% ��Jo�o#5GY  o}���o��������m   �iN�`�r����������̏ޏ����   $�,�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�bϸtφ��  
�`(�  �B�( 	 ���Ϻ������ �8�&�H�J�\ߒ߀�жߤ��ߠ�4� �n�1�C�g�y� �������c����� �V�3�E�W�i�{��� ���������� /AS��w���� ����`r Oas����� ��8/'/9/�]/ o/�/�/�/�/��/�/ �/F/#?5?G?Y?k?}? �/�/�?�?�??�?O O1OCOUO�?yO�O�O �?�O�O�O�O	__bO ?_Q_c_�O�_�_�_�_ �_�_(_:_o)o;o�_ _oqo�o�o�o�o o�o �oHo%7I[m �o����� �!�3�E���{��� ���ÏՏ����� d�A�S�e��������� ��џ�*���+�r� O�a�s����������@ ˢد���ˣ�ҧ����)fr�h:\tpgl\�robots\r�2000ic6�_�165f.xml ��`�r���������̿0޿������3� E�W�i�{ύϟϱ��� �������
�/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�9�K�]�o����� �������������# 5GYk}��� ��� �1C Ugy����� ���/-/?/Q/c/ u/�/�/�/�/�/�/�.:�K� ү ��<< �?��+6?�/.?P?~?d? �?�?�?�?�?�?�?O 2OO:OhONO`O�O�O�O�O�O���$TP�GL_OUTPU�T ���� 0U3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�oU0���@2345678901�o, >PXs���o�� ���q��!�3�E�W��z}a������� ��яi�{���+�=� O�a���o�������͟ ߟw���'�9�K�]� ���������ɯۯ� ����#�5�G�Y�k�� y�����ſ׿鿁��� �1�C�U�g�y�χ� ���������Ϗ��-� ?�Q�c�u��߽߫� ���������;�M� _�q���������������A}17�I� [�m������@?�����: ( 	 �o��1UC yg������ �	?-Ouc �������� /;/)/_/�f�0-6 g/�/�-�/�/�/�/? ?�j�/F?X?�/d?�? h?z?�?�?4?�?O�? �?BOTO.OxO�O�?rO �OZO�O�O_�O,_>_ �O&_t_�_ _�_�_�_ �_�_P_b_(o:o�_Bo poJo\o�o�oo�o�o �o�o$�oZl�o t�<�����  �~�V�h������ x���ԏ2���
���� @�R�,�>�������� Пj�ܟ����<�N� ��R����p���̯�� ��`��8�ү$�n� ��Z����������� ��"�4��@�j�ȿڿ �ϲ�LϺ�������� 0ߎ�T�f� �Rߜ�v��������v"�$TP�OFF_LIM �{ ��w!������N_SV� � ���P_M�ON s%�����2����S�TRTCHK �s%�4��VT?COMPAT*����VWVAR �J���.� R�� ���]����_DEFPROG� %y�%F�GF _1���_DISPLAY
��y��INST_M�SK  q� ~[�INUSER���a�LCK��z�QU?ICKMEN��a�oSCRE��s%~��tpsca���� 	�' _+	S�T���RACE_�CFG J�����	��
?�~rHNL 2.�S ��� ����� $6HZtI�TEM 2�� �%$1234?567890��  =<�����  !��� �:/��[/�/�/ ��//+/�/O/?s/ ?E?�/�/�/�/�/? }?'?�?�?Oo?/O�? �?�?1O�?�O�O�O#O �OGOYOkO�O=_�Oa_ s_�O_�O_�_1_�_ U_o'o�_=o�_o�o �_�o	o�o�o�oQo�o uo�o�o�oi�� �);M��� C�U��a������ ӏ7���	�m������ l�Ǐ��돗���C�3� E�W�q�{�����K�q� ��矧���/���S� ��%�7���C���ѯ� g����ٿ�O���s� ��Nϩ�i�Ϳ�ϟ�� ��'�y��]�߁�-� S�e���q�����ߋ� 5�����}�=�߳� ��I�a��߻���1��� U�g�0���K���o���@���	����pS|�����  �e�� �@7�
� MsZ�
�UD1:\������R_GRP 1��� 	 @@���!E3iW�y���c�����?�  /+/9/'/]/ K/�/o/�/�/�/�/�/ �/�/#??G?5?W?}?�	���?�?��SC�B 2  ��?OO%O7OIO[O�mOO��UTORIAL ��O���V_CONFIG �=��)_�MOUTPUT� 	P��5_y_�_�_�_�_�_ �_�_	oo-o?oQoQ f_yo�o�o�o�o�o�o �o	-?Qbou �������� �)�;�M�^q����� ����ˏݏ���%� 7�I�[�l�������� ǟٟ����!�3�E� W�h�{�������ïկ �����/�A�S�d� w���������ѿ��� ��+�=�O�a�r��� �ϩϻ��������� '�9�K�]�nρߓߥ� �����������#�5� G�Y�j�}������ ��������1�C�U� g�_Ud_�������� ����#5GYk }p������ 1CUgy� ������	// -/?/Q/c/u/�/��/ �/�/�/�/??)?;? M?_?q?�?�/�?�?�? �?�?OO%O7OIO[O mOO�?�O�O�O�O�O �O_!_3_E_W_i_{_ �_�O�_�_�_�_�_o o/oAoSoeowo�o�_ �o�o�o�o�o+ =Oas��o�� �����'�9�K� ]�o��������ɏۏ ����#�5�G�Y�k��}���r���� ��������럎��!� 3�E�W�i�{������� ïկ篚���/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�o߁� �ߥ߷���������� #�5�G�Y�k�}��� ������������1� C�U�g�y��������� �������-?Q cu������ �);M_q �������/ %/7/I/[/m//�/ �/�/�/�/�/�//!? 3?E?W?i?{?�?�?�?��?�?�?�?K�$T�X_SCREEN� 1���}�OLO^OpO�O�O�O:O��9O �O�O
__._@_�O�O v_�_�_�_�_�_G_�_ k_o*o<oNo`oro�_ �oo�o�o�o�o �o�oJ\n��� �?���"�4� F��j��������ď ֏�_�q��0�B�T� f�x�����ҟ��������>��$U�ALRM_MSG� ?(I�5@  6�:p�������ׯʯ ��� ��$�U�H�y��l���Q�SEV  �_�϶O�EC�FG (E�2A  5@� � A��   B�4
 ��3(E2� D�V�h�zόϞϰ����������۱GRP �2� 06	� �>�Q�I_B�BL_NOTE � �T�G�l2-@1�~Q�DEFPRO[�=%_� (%���� 0���������'�� K�6�\��l������G�FKEYDAT�A 1!(I(�ps ��6 �π-�?�|��f�x�R�,(���4�������� ��.R9v� o������ *<#`G�k�0�������/ '/9/K/]/o/2/�/ �/�/�/�/�/�/?(? :?L?^?p?�/�?�?�? �?�?�? O�?$O6OHO ZOlO~OO�O�O�O�O �O�O�O _2_D_V_h_ z_�__�_�_�_�_�_ 
o�_.o@oRodovo�o o�o�o�o�o�o �o<N`r��% �������8� J�\�n�������3�ȏ ڏ����"��F�X� j�|�������ğ֟� ����0���T�f�x� ������=�ү���� �,���P�b�t����� ����K�����(� :�ɿ^�pςϔϦϸ� G����� ��$�6�H� ��l�~ߐߢߴ���U� ����� �2�D���h� z��������c��� 
��.�@�R���v��� ��������_����*<N`7�f}�;�����@������,� �<#`rY� }�����/&/ /J/1/n/�/g/�/�/ �/�/�/�/�/"?	?F? X?7�|?�?�?�?�?�? ���?OO0OBOTOfO �?�O�O�O�O�O�OsO __,_>_P_b_�O�_ �_�_�_�_�_�_�_o (o:oLo^opo�_�o�o �o�o�o�o}o$6 HZl~��� ���� �2�D�V� h�z�	�����ԏ� ��
���.�@�R�d�v� �������П���� ��*�<�N�`�r����� m?��̯ޯ���� 8�J�\�n�������3� ȿڿ����"ϱ�F� X�j�|ώϠ�/����� ������0߿�T�f� xߊߜ߮�=������� ��,��P�b�t�� ����K������� (�:���^�p������� ��G����� $6 H��l~���� U�� 2D� hz����������������/#-�E/W/1&,C?�/;?�/�/�/ �/�/?�/*?<?#?`? G?�?�?}?�?�?�?�? �?O�?8OO\OnOUO �OyO�O�O���O�O_ "_4_F_Uj_|_�_�_ �_�_�_e_�_oo0o BoTo�_xo�o�o�o�o �oao�o,>P b�o������ o��(�:�L�^�� ��������ʏ܏�}� �$�6�H�Z�l����� ����Ɵ؟�y�� � 2�D�V�h�z�	����� ¯ԯ������.�@� R�d�v��������п �����O*�<�N�`� rτϋ��Ϻ������� �ߣ�8�J�\�n߀� ��!߶���������� ��4�F�X�j�|��� /������������� B�T�f�x�����+��� ������,��P bt���9�� �(�L^p ����G�� / /$/6/�Z/l/~/�/ �/�/C/�/�/�/? ?h2?D?�F;�����o?�?�=k?�?�?�6,�O�?�O OO@ORO9OvO]O�O �O�O�O�O�O_�O*_ _N_`_G_�_k_�_�_ �_�_�_o�_&o8o� \ono�o�o�o�o�/�o �o�o"4F�oj |����S�� ��0�B��f�x��� ������ҏa����� ,�>�P�ߏt������� ��Ο]����(�:� L�^�ퟂ�������ʯ ܯk� ��$�6�H�Z� �~�������ƿؿ� y�� �2�D�V�h��� �Ϟϰ�������u�
� �.�@�R�d�v�Mo�� �߾����������*� <�N�`�r����� ���������&�8�J� \�n������������ ������4FXj |������ �0BTfx� �+����// �>/P/b/t/�/�/'/ �/�/�/�/??(?�/ L?^?p?�?�?�?5?�? �?�? OO$O�?HOZO@lO~O�O�O�O���K���������O�O]�O%_7_V, #oh_o�_s_�_�_�_ �_�_
ooo@o'odo vo]o�o�o�o�o�o�o �o�o<N5rY ��������� &�5OJ�\�n������� ��E�ڏ����"�4� ÏX�j�|�������A� ֟�����0�B�џ f�x���������O�� ����,�>�ͯb�t� ��������ο]��� �(�:�L�ۿpςϔ� �ϸ���Y��� ��$� 6�H�Z���~ߐߢߴ� ����g���� �2�D� V���z�������� ��
��.�@�R�d� k�������������� ��*<N`r ������ &8J\n�� ������"/4/ F/X/j/|//�/�/�/ �/�/�/?�/0?B?T? f?x?�??�?�?�?�? �?O�?,O>OPObOtO �O�O'O�O�O�O�O_ _�O:_L_^_p_�_�_ #_�_�_�_�_ oo$o���&k������OoaosmKo�o�o�f,��o��o�o  2V=z�s �����
��.� @�'�d�K���o����� ���ɏ����<�N� `�r������_��̟ޟ ���&���J�\�n� ������3�ȯگ��� �"���F�X�j�|��� ����A�ֿ����� 0Ͽ�T�f�xϊϜϮ� =���������,�>� ��b�t߆ߘߪ߼�K� ������(�:���^� p�������Y���  ��$�6�H���l�~� ��������U�����  2DV-�z�� ������
. @Rd����� ��q//*/</N/ `/��/�/�/�/�/�/ �//?&?8?J?\?n? �/�?�?�?�?�?�?{? O"O4OFOXOjO|OO �O�O�O�O�O�O�O_ 0_B_T_f_x__�_�_ �_�_�_�_o�_,o>o Poboto�oo�o�o�o �o�o�o(:L^�p��k �{�>k ����� �}����v,�H� ��l�S�������Ə�� ���� ��D�V�=� z�a�������ԟ���� ߟ�.��R�9�v��� g����Я���� *�<�N�`�r�����%� ��̿޿��ϣ�8� J�\�nπϒ�!϶��� �������"߱�F�X� j�|ߎߠ�/������� �����B�T�f�x� ����=�������� �,���P�b�t����� ��9�������( :��^p���� G�� $6� Zl~������ ��/ /2/D/Kh/ z/�/�/�/�/�/c/�/ 
??.?@?R?�/v?�? �?�?�?�?_?�?OO *O<ONO`O�?�O�O�O �O�O�OmO__&_8_ J_\_�O�_�_�_�_�_ �_�_{_o"o4oFoXo jo�_�o�o�o�o�o�o wo0BTfx ������� �,�>�P�b�t���������Ώ������������/�A�S�+�u���a�,s���k�ܟß �� ��6��Z�l�S���w� ��Ư���ѯ� �� D�+�h�O�������¿ �������.�@�R� d�vυ��ϬϾ����� ��ߕ�*�<�N�`�r� ��ߨߺ�������� ��&�8�J�\�n��� !������������� 4�F�X�j�|������ ����������B Tfx��+�� ���>Pb t���9��� //(/�L/^/p/�/ �/�/5/�/�/�/ ?? $?6?�Z?l?~?�?�? �?�/�?�?�?O O2O DO�?hOzO�O�O�O�O QO�O�O
__._@_�O d_v_�_�_�_�_�___ �_oo*o<oNo�_ro �o�o�o�o�o[o�o &8J\�o�� ����i��"� 4�F�X��|������� ď֏�w���0�B� T�f�����������ҟ �s���,�>�P�b��t�K0v��K0�������í�����Ѧ,�(�ۿL� 3�p���i�����ʿܿ ÿ ��$�6��Z�A� ~ϐ�wϴϛ��Ͽ��� ���2��V�h�G?�� �߰���������
�� .�@�R�d�v���� ����������*�<� N�`�r���������� ������&8J\ n������ ��"4FXj| ������/ �0/B/T/f/x/�// �/�/�/�/�/??�/ >?P?b?t?�?�?'?�? �?�?�?OO�?:OLO ^OpO�O�O�O}��O�O �O __$_+OH_Z_l_ ~_�_�_�_C_�_�_�_ o o2o�_Vohozo�o �o�o?o�o�o�o
 .@�odv��� �M����*�<� �`�r���������̏ [�����&�8�J�ُ n���������ȟW�� ���"�4�F�X��|� ������į֯e���� �0�B�T��x��������ҿ��$UI�_INUSER � ������  ���_MENHI�ST 1"��  ( ����(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1$ϗϩϜ���π� _�q�936���+�=�O��� f�xߊߜ߮�����a� ����,�>�P���t� �������]���� �(�:�L�^������ ��������k� $6HZj���Y��� �������� &8J\n��� ����{�"/4/ F/X/j/|//�/�/�/ �/�/�/�/?0?B?T? f?x???�?�?�?�? �?O�?,O>OPObOtO �Oq��O�O�O�O_ _O:_L_^_p_�_�_ #_�_�_�_�_ oo$o �_HoZolo~o�o�o1o �o�o�o�o �oD Vhz���?� ��
��.��R�d� v��������O�O�� ��*�<�?�`�r��� ������I�ޟ��� &�8�J�ٟn������� ��ȯW�����"�4� F�կj�|�������Ŀ ֿe�����0�B�T� �xϊϜϮ����Ͻ� Ϗ��,�>�P�b�e� �ߘߪ߼�����o߁� �(�:�L�^�p��ߔ� ���������}��$� 6�H�Z�l�������� ���������� 2D Vhz	�����������$UI�_PANEDAT�A 1$����.  	��}  frh�/cgtp/fl�exdev.st�m?_width�=0&_heig�ht=10^Oi�ce=TP&_l�ines=15&�_columns�=4^font=�24&_page?=wholeO
~��)  rim��  ?��/#/ 5/G/�Y/}/d/�/�/ �/�/�/�/�/?1??�U?<?y?�?r?�?��� ���2��?�? OO1OCO�?gO�yO �O�O�O�O�O�O^O_ _?_&_Q_u_\_�_�_ �_�_�_�_�_o)ooMo�<nf0�O�o�o �o�o�o�o=o�O2 DVhz��o�� ���
���@�'� d�K������������ �goyo*�<�N�`�r� ��׏��̟ޟ�� �&�8���\�C���g� ������گ������� 4��X�j�Q����� Ŀֿ�����q�B� T�ǟxϊϜϮ����� 9������,��P�7� t߆�mߪߑ������� ���(��k�p�� ���������a�� $�6�H�Z�l������ ������������  D+hza��� �G�Y�
.@R d������� �//</#/`/G/ �/�/}/�/�/�/�/�/ ?�/8?J?1?n?�� �?�?�?�?�?�?Q?"O 4O�XOjO|O�O�O�O O�O�O�O_�O0__ T_f_M_�_q_�_�_�_`�_�_o{?�?}�o@Rodovo�o�o�o)@o �oDE�o�o!3E W�o{b���� ����/��S�:��w���p���=H�3�;��$UI_POST�YPE  �5�� 	 ����߂QUICK�MEN  ������RESTO�RE 1%�5�  ����FB������FBm ��ޟ���&�ɟJ� \�n�����5���ȯگ �������/���j� |�������U�ֿ��� ��0�ӿT�f�xϊ� ��G��ϻ���?��� ,�>�P���t߆ߘߪ� ��_�������(��� ��G�Y���}����� ������$�6�H�Z� ��~���������q��� ����i�2DVhz ��������.@Rd�SC�RE.�?3��u1sc�uU2�3�4�5��6�7�8�|T;AT�� B��5׊USER����T��ks�:$4�:$5:$6:$7:$8�:!߀NDO_CFG &�)`(a߀�PD�)�None ߀� _INFO 1�'�5� @�0% j�/=H�/?�/4?F? )?j?|?_?�?�?�?�?��?�?O�?0O��!O�FFSET *��!=Ox��O �O�O�O�O�O�O__ #_mO'_t_k_}_�_�_ �_�_�_�_�_E[C�Gm�5ojo
Zo�oIHUFRAME  ��&�!RTOL_�ABRT�oMC�bE�NB�o�hGRP �1+s�?�Cz  A�*s(q�!(: L^p���{�f-��U�h�!�kMSK � �e�!�kN�a�r� �%o8� �VC�MRr21_K��y	� B�1: SC130EF2 *����e�DX��$�t�5��!?��p@�pp:�p�<� ~o����'�T�y�O��|���uA��h��� B���ԑؕ`���@� ��A�,�e�P���t� �����������+��ޟO�a�J�ISIO�NTMOU�`�t�%�x�t"2SﳸS� q FR:\z��\� A\f� �߀ MC��LO�Gƿ   UD�1��EX�'� B@ �� -���'�K���O�s�� � n6  ����*��t��`���  =���������}߸TRAINϸ����|`  d�Qp�ə�U�3_M(� ��E��E�S�e�w߉� �߭�����������h+�=�r�_�RE���4y�J�LEXEr��5_K�!1-eh��VMPHAS��%�#АK�RTD�_FILTER �26_K �GU� �0�B�T�f�x����� ������BZ�' 9K]o���H��SHIFT�r17_K
 <:�&�� ��=&sJ \��������'/�/]/4/	L�IVE/SNAP�Cvsfliv\��o/�z� Y@yU� �"menu�/��/G/??�"���8X�	��MO��9���ĵp�$WAIT?DINEND���x�~4O�p��7���?S��?�9TIM�u���<G�?M�?6K�?�J�?JO�8REL�E���o{4����~1_ACT� �H ��B± :� ?F_�f�B�RDIS� �o�$�XVR��;���_$ZABCs<�� ,|h2N_�mZ[IP��=����o(o:o�ZMPCF�_G 1>{ A0��o�oRgs?y�q� ���o;�7<�� �o
 ��o@�gԁ2�]C -�Qs����Х�Հ)�#�5�K�Y����P[`��@�_�S�P_YLIND �Ack� ��,(  *���9����B�)� �x�����ޏ ��.��ʟܟ�\�=� O�a����� �������߯Ư4��'��[�c29BcgQ �xor� ���������Ͽ�yb�����w��A4���S�PHERE 2Cč�y�U�ɯNϋ�r� ����
�����s�ߺ� ��Q�8�u�\��ϫ߽� ����f�����M�`��q���PZZ�F ��F